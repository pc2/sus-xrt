// THIS IS A GENERATED FILE (Generated at 2025-11-26T15:04:41+01:00)
// This file was generated with SUS Compiler 0.3.6 () built at 2025-11-13_15:28:01 
// all_benchmarks #()
module all_benchmarks(
	input clk
);

benchmark_burst_read_AXI_WIDTH_32 burst32(
	.aclk(clk),
	.aresetn(),
	.s_axi_control_awaddr(),
	.s_axi_control_awvalid(),
	.s_axi_control_awready(),
	.s_axi_control_wdata(),
	.s_axi_control_wstrb(),
	.s_axi_control_wvalid(),
	.s_axi_control_wready(),
	.s_axi_control_bresp(),
	.s_axi_control_bvalid(),
	.s_axi_control_bready(),
	.s_axi_control_araddr(),
	.s_axi_control_arvalid(),
	.s_axi_control_arready(),
	.s_axi_control_rdata(),
	.s_axi_control_rresp(),
	.s_axi_control_rvalid(),
	.s_axi_control_rready(),
	.m_axi_awvalid(),
	.m_axi_awready(),
	.m_axi_awaddr(),
	.m_axi_awlen(),
	.m_axi_awburst(),
	.m_axi_awcache(),
	.m_axi_wvalid(),
	.m_axi_wready(),
	.m_axi_wdata(),
	.m_axi_wstrb(),
	.m_axi_wlast(),
	.m_axi_bvalid(),
	.m_axi_bready(),
	.m_axi_bresp(),
	.m_axi_arvalid(),
	.m_axi_arready(),
	.m_axi_araddr(),
	.m_axi_arlen(),
	.m_axi_arsize(),
	.m_axi_arburst(),
	.m_axi_rvalid(),
	.m_axi_rready(),
	.m_axi_rdata(),
	.m_axi_rresp(),
	.m_axi_rlast(),
	.m_axi_arprot(),
	.m_axi_arcache(),
	.m_axi_arqos(),
	.m_axi_arlock(),
	.m_axi_arregion()
);
benchmark_burst_read_AXI_WIDTH_64 burst64(
	.aclk(clk),
	.aresetn(),
	.s_axi_control_awaddr(),
	.s_axi_control_awvalid(),
	.s_axi_control_awready(),
	.s_axi_control_wdata(),
	.s_axi_control_wstrb(),
	.s_axi_control_wvalid(),
	.s_axi_control_wready(),
	.s_axi_control_bresp(),
	.s_axi_control_bvalid(),
	.s_axi_control_bready(),
	.s_axi_control_araddr(),
	.s_axi_control_arvalid(),
	.s_axi_control_arready(),
	.s_axi_control_rdata(),
	.s_axi_control_rresp(),
	.s_axi_control_rvalid(),
	.s_axi_control_rready(),
	.m_axi_awvalid(),
	.m_axi_awready(),
	.m_axi_awaddr(),
	.m_axi_awlen(),
	.m_axi_awburst(),
	.m_axi_awcache(),
	.m_axi_wvalid(),
	.m_axi_wready(),
	.m_axi_wdata(),
	.m_axi_wstrb(),
	.m_axi_wlast(),
	.m_axi_bvalid(),
	.m_axi_bready(),
	.m_axi_bresp(),
	.m_axi_arvalid(),
	.m_axi_arready(),
	.m_axi_araddr(),
	.m_axi_arlen(),
	.m_axi_arsize(),
	.m_axi_arburst(),
	.m_axi_rvalid(),
	.m_axi_rready(),
	.m_axi_rdata(),
	.m_axi_rresp(),
	.m_axi_rlast(),
	.m_axi_arprot(),
	.m_axi_arcache(),
	.m_axi_arqos(),
	.m_axi_arlock(),
	.m_axi_arregion()
);
benchmark_burst_read_AXI_WIDTH_128 burst128(
	.aclk(clk),
	.aresetn(),
	.s_axi_control_awaddr(),
	.s_axi_control_awvalid(),
	.s_axi_control_awready(),
	.s_axi_control_wdata(),
	.s_axi_control_wstrb(),
	.s_axi_control_wvalid(),
	.s_axi_control_wready(),
	.s_axi_control_bresp(),
	.s_axi_control_bvalid(),
	.s_axi_control_bready(),
	.s_axi_control_araddr(),
	.s_axi_control_arvalid(),
	.s_axi_control_arready(),
	.s_axi_control_rdata(),
	.s_axi_control_rresp(),
	.s_axi_control_rvalid(),
	.s_axi_control_rready(),
	.m_axi_awvalid(),
	.m_axi_awready(),
	.m_axi_awaddr(),
	.m_axi_awlen(),
	.m_axi_awburst(),
	.m_axi_awcache(),
	.m_axi_wvalid(),
	.m_axi_wready(),
	.m_axi_wdata(),
	.m_axi_wstrb(),
	.m_axi_wlast(),
	.m_axi_bvalid(),
	.m_axi_bready(),
	.m_axi_bresp(),
	.m_axi_arvalid(),
	.m_axi_arready(),
	.m_axi_araddr(),
	.m_axi_arlen(),
	.m_axi_arsize(),
	.m_axi_arburst(),
	.m_axi_rvalid(),
	.m_axi_rready(),
	.m_axi_rdata(),
	.m_axi_rresp(),
	.m_axi_rlast(),
	.m_axi_arprot(),
	.m_axi_arcache(),
	.m_axi_arqos(),
	.m_axi_arlock(),
	.m_axi_arregion()
);
benchmark_burst_read_AXI_WIDTH_256 burst256(
	.aclk(clk),
	.aresetn(),
	.s_axi_control_awaddr(),
	.s_axi_control_awvalid(),
	.s_axi_control_awready(),
	.s_axi_control_wdata(),
	.s_axi_control_wstrb(),
	.s_axi_control_wvalid(),
	.s_axi_control_wready(),
	.s_axi_control_bresp(),
	.s_axi_control_bvalid(),
	.s_axi_control_bready(),
	.s_axi_control_araddr(),
	.s_axi_control_arvalid(),
	.s_axi_control_arready(),
	.s_axi_control_rdata(),
	.s_axi_control_rresp(),
	.s_axi_control_rvalid(),
	.s_axi_control_rready(),
	.m_axi_awvalid(),
	.m_axi_awready(),
	.m_axi_awaddr(),
	.m_axi_awlen(),
	.m_axi_awburst(),
	.m_axi_awcache(),
	.m_axi_wvalid(),
	.m_axi_wready(),
	.m_axi_wdata(),
	.m_axi_wstrb(),
	.m_axi_wlast(),
	.m_axi_bvalid(),
	.m_axi_bready(),
	.m_axi_bresp(),
	.m_axi_arvalid(),
	.m_axi_arready(),
	.m_axi_araddr(),
	.m_axi_arlen(),
	.m_axi_arsize(),
	.m_axi_arburst(),
	.m_axi_rvalid(),
	.m_axi_rready(),
	.m_axi_rdata(),
	.m_axi_rresp(),
	.m_axi_rlast(),
	.m_axi_arprot(),
	.m_axi_arcache(),
	.m_axi_arqos(),
	.m_axi_arlock(),
	.m_axi_arregion()
);
benchmark_burst_read_AXI_WIDTH_512 burst512(
	.aclk(clk),
	.aresetn(),
	.s_axi_control_awaddr(),
	.s_axi_control_awvalid(),
	.s_axi_control_awready(),
	.s_axi_control_wdata(),
	.s_axi_control_wstrb(),
	.s_axi_control_wvalid(),
	.s_axi_control_wready(),
	.s_axi_control_bresp(),
	.s_axi_control_bvalid(),
	.s_axi_control_bready(),
	.s_axi_control_araddr(),
	.s_axi_control_arvalid(),
	.s_axi_control_arready(),
	.s_axi_control_rdata(),
	.s_axi_control_rresp(),
	.s_axi_control_rvalid(),
	.s_axi_control_rready(),
	.m_axi_awvalid(),
	.m_axi_awready(),
	.m_axi_awaddr(),
	.m_axi_awlen(),
	.m_axi_awburst(),
	.m_axi_awcache(),
	.m_axi_wvalid(),
	.m_axi_wready(),
	.m_axi_wdata(),
	.m_axi_wstrb(),
	.m_axi_wlast(),
	.m_axi_bvalid(),
	.m_axi_bready(),
	.m_axi_bresp(),
	.m_axi_arvalid(),
	.m_axi_arready(),
	.m_axi_araddr(),
	.m_axi_arlen(),
	.m_axi_arsize(),
	.m_axi_arburst(),
	.m_axi_rvalid(),
	.m_axi_rready(),
	.m_axi_rdata(),
	.m_axi_rresp(),
	.m_axi_rlast(),
	.m_axi_arprot(),
	.m_axi_arcache(),
	.m_axi_arqos(),
	.m_axi_arlock(),
	.m_axi_arregion()
);
axi_realigning_burst_reader_T_type_bool_32_17_AXI_WIDTH_512_ADDR_ALIGN_4_COUNT_TO_65536_ATO_18446744073709551616 reader_for_testbench(
	.aclk(clk),
	.aresetn(),
	.arvalid(),
	.arready(),
	.araddr(),
	.arlen(),
	.arsize(),
	.arburst(),
	.arprot(),
	.arcache(),
	.arqos(),
	.arlock(),
	.arregion(),
	.rvalid(),
	.rready(),
	.rdata(),
	.rresp(),
	.rlast(),
	.max_in_flight(),
	.may_request_new_burst(),
	.request_new_burst(),
	.start_addr(),
	.count(),
	.is_ready_to_receive_lots_of_data(),
	.value_valid(),
	.value(),
	.last()
);
endmodule

// benchmark_burst_read #(AXI_WIDTH: 512)
module benchmark_burst_read_AXI_WIDTH_512(
	input aclk,
	input wire aresetn,
	input wire[11:0] s_axi_control_awaddr,
	input wire s_axi_control_awvalid,
	output /*mux_wire*/ logic s_axi_control_awready,
	input wire[31:0] s_axi_control_wdata,
	input wire[3:0] s_axi_control_wstrb,
	input wire s_axi_control_wvalid,
	output /*mux_wire*/ logic s_axi_control_wready,
	output /*mux_wire*/ logic[1:0] s_axi_control_bresp,
	output /*mux_wire*/ logic s_axi_control_bvalid,
	input wire s_axi_control_bready,
	input wire[11:0] s_axi_control_araddr,
	input wire s_axi_control_arvalid,
	output /*mux_wire*/ logic s_axi_control_arready,
	output /*mux_wire*/ logic[31:0] s_axi_control_rdata,
	output /*mux_wire*/ logic[1:0] s_axi_control_rresp,
	output /*mux_wire*/ logic s_axi_control_rvalid,
	input wire s_axi_control_rready,
	output /*mux_wire*/ logic m_axi_awvalid,
	input wire m_axi_awready,
	output /*mux_wire*/ logic[63:0] m_axi_awaddr,
	output /*mux_wire*/ logic[7:0] m_axi_awlen,
	output /*mux_wire*/ logic[1:0] m_axi_awburst,
	output /*mux_wire*/ logic[3:0] m_axi_awcache,
	output /*mux_wire*/ logic m_axi_wvalid,
	input wire m_axi_wready,
	output /*mux_wire*/ logic[511:0] m_axi_wdata,
	output /*mux_wire*/ logic[63:0] m_axi_wstrb,
	output /*mux_wire*/ logic m_axi_wlast,
	input wire m_axi_bvalid,
	output /*mux_wire*/ logic m_axi_bready,
	input wire[1:0] m_axi_bresp,
	output /*mux_wire*/ logic m_axi_arvalid,
	input wire m_axi_arready,
	output /*mux_wire*/ logic[63:0] m_axi_araddr,
	output /*mux_wire*/ logic[7:0] m_axi_arlen,
	output /*mux_wire*/ logic[2:0] m_axi_arsize,
	output /*mux_wire*/ logic[1:0] m_axi_arburst,
	input wire m_axi_rvalid,
	output /*mux_wire*/ logic m_axi_rready,
	input wire[511:0] m_axi_rdata,
	input wire[1:0] m_axi_rresp,
	input wire m_axi_rlast,
	output /*mux_wire*/ logic[2:0] m_axi_arprot,
	output /*mux_wire*/ logic[3:0] m_axi_arcache,
	output /*mux_wire*/ logic[3:0] m_axi_arqos,
	output /*mux_wire*/ logic m_axi_arlock,
	output /*mux_wire*/ logic[3:0] m_axi_arregion
);

genvar _g0;
/*mux_wire*/ logic _ctrl_aresetn;
wire _ctrl_awready;
wire _ctrl_wready;
wire[1:0] _ctrl_bresp;
wire _ctrl_bvalid;
wire _ctrl_arready;
wire[31:0] _ctrl_rdata;
wire[1:0] _ctrl_rresp;
wire _ctrl_rvalid;
/*mux_wire*/ logic[11:0] _ctrl_awaddr;
/*mux_wire*/ logic _ctrl_awvalid;
/*mux_wire*/ logic[31:0] _ctrl_wdata;
/*mux_wire*/ logic[3:0] _ctrl_wstrb;
/*mux_wire*/ logic _ctrl_wvalid;
/*mux_wire*/ logic _ctrl_bready;
/*mux_wire*/ logic[11:0] _ctrl_araddr;
/*mux_wire*/ logic _ctrl_arvalid;
/*mux_wire*/ logic _ctrl_rready;
/*mux_wire*/ logic _reader_aresetn;
/*mux_wire*/ logic _writer_aresetn;
wire _writer_awvalid;
wire[63:0] _writer_awaddr;
wire[7:0] _writer_awlen;
wire[1:0] _writer_awburst;
wire[3:0] _writer_awcache;
wire _writer_wvalid;
wire[511:0] _writer_wdata;
wire[63:0] _writer_wstrb;
wire _writer_wlast;
wire _writer_bready;
/*mux_wire*/ logic _writer_awready;
/*mux_wire*/ logic _writer_wready;
/*mux_wire*/ logic _writer_bvalid;
/*mux_wire*/ logic[1:0] _writer_bresp;
wire _reader_arvalid;
wire[63:0] _reader_araddr;
wire[7:0] _reader_arlen;
wire[2:0] _reader_arsize;
wire[1:0] _reader_arburst;
wire _reader_rready;
/*mux_wire*/ logic _reader_arready;
/*mux_wire*/ logic _reader_rvalid;
/*mux_wire*/ logic[511:0] _reader_rdata;
/*mux_wire*/ logic[1:0] _reader_rresp;
/*mux_wire*/ logic _reader_rlast;
/*mux_wire*/ logic[63:0] addr_a_bits;
wire[31:0] _ctrl_input_regs[3:0];
wire[31:0] _46 = _ctrl_input_regs[0];
wire[31:0] _47 = _ctrl_input_regs[1];
/*mux_wire*/ logic[63:0] start_addr;
/*mux_wire*/ logic[63:0] _BitsToUInt_bits;
wire[63:0] _BitsToUInt_value;
/*mux_wire*/ logic[31:0] num_to_transfer;
wire[31:0] _49 = _ctrl_input_regs[2];
/*mux_wire*/ logic[31:0] _BitsToUInt_2_bits;
wire[31:0] _BitsToUInt_2_value;
/*mux_wire*/ logic[31:0] _IntNarrow_in;
wire[31:0] _IntNarrow_out;
/*mux_wire*/ logic[31:0] config_bits;
wire[31:0] _50 = _ctrl_input_regs[3];
wire[2:0] _51;
generate
for(_g0 = 0; _g0 < 3; _g0 = _g0 + 1) begin
assign _51[_g0] = config_bits[5 + _g0];
end
endgenerate
wire[3:0] _52;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _52[_g0] = config_bits[8 + _g0];
end
endgenerate
wire[3:0] _53;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _53[_g0] = config_bits[12 + _g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_3_bits;
wire[3:0] _BitsToUInt_3_value;
wire _54 = config_bits[16];
wire[3:0] _55;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _55[_g0] = config_bits[17 + _g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_4_bits;
wire[3:0] _BitsToUInt_4_value;
wire[10:0] _56;
generate
for(_g0 = 0; _g0 < 11; _g0 = _g0 + 1) begin
assign _56[_g0] = config_bits[21 + _g0];
end
endgenerate
/*mux_wire*/ logic[10:0] _BitsToUInt_5_bits;
wire[10:0] _BitsToUInt_5_value;
/*mux_wire*/ logic[10:0] _reader_max_in_flight;
/*state*/ logic[63:0] cycles_since_reset;
wire[64:0] _59;
assign _59 = cycles_since_reset + 1'd1;
wire[63:0] _60;
assign _60 = _59; // == mod 18446744073709551616 (target is 64 bits wide)
/*mux_wire*/ logic[63:0] cycles_since_reset_bits;
/*mux_wire*/ logic[63:0] _UIntToBits_value;
wire[63:0] _UIntToBits_bits;
/*latency*/ logic[63:0] __UIntToBits_bits_D1; always_ff @(posedge aclk) begin __UIntToBits_bits_D1 <= _UIntToBits_bits; end
/*latency*/ logic[63:0] __UIntToBits_bits_D2; always_ff @(posedge aclk) begin __UIntToBits_bits_D2 <= __UIntToBits_bits_D1; end
/*latency*/ logic[63:0] __UIntToBits_bits_D3; always_ff @(posedge aclk) begin __UIntToBits_bits_D3 <= __UIntToBits_bits_D2; end
/*state*/ logic[63:0] cycles_since_reset_at_start;
/*state*/ logic running;
/*state*/ logic[31:0] num_cycles_running;
/*state*/ logic[31:0] hash;
wire _ctrl_start;
/*latency*/ logic __ctrl_start_D1; always_ff @(posedge aclk) begin __ctrl_start_D1 <= _ctrl_start; end
/*latency*/ logic __ctrl_start_D2; always_ff @(posedge aclk) begin __ctrl_start_D2 <= __ctrl_start_D1; end
/*latency*/ logic __ctrl_start_D3; always_ff @(posedge aclk) begin __ctrl_start_D3 <= __ctrl_start_D2; end
/*mux_wire*/ logic _reader_request_new_burst;
/*mux_wire*/ logic[63:0] _reader_start_addr;
/*mux_wire*/ logic[31:0] _reader_count;
localparam[31:0] _67 = 32'b00000000000000000000000000000000;
wire[32:0] _72;
assign _72 = num_cycles_running + 1'd1;
wire[31:0] _73;
assign _73 = _72; // == mod 4294967296 (target is 32 bits wide)
/*mux_wire*/ logic _reader_is_ready_to_receive_lots_of_data;
wire _reader_value_valid;
/*latency*/ logic __reader_value_valid_D1; always_ff @(posedge aclk) begin __reader_value_valid_D1 <= _reader_value_valid; end
/*latency*/ logic __reader_value_valid_D2; always_ff @(posedge aclk) begin __reader_value_valid_D2 <= __reader_value_valid_D1; end
/*latency*/ logic __reader_value_valid_D3; always_ff @(posedge aclk) begin __reader_value_valid_D3 <= __reader_value_valid_D2; end
wire[31:0] _reader_value[15:0];
wire _reader_last;
/*mux_wire*/ logic[31:0] value[15:0];
/*mux_wire*/ logic last;
/*latency*/ logic _last_D1; always_ff @(posedge aclk) begin _last_D1 <= last; end
/*latency*/ logic _last_D2; always_ff @(posedge aclk) begin _last_D2 <= _last_D1; end
/*latency*/ logic _last_D3; always_ff @(posedge aclk) begin _last_D3 <= _last_D2; end
/*mux_wire*/ logic[31:0] new_hash_contrib;
wire[15:0] _74;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _74[_g0] = value[_g0][0];
end
endgenerate
wire _75;
assign _75 = ^_74;
/*latency*/ logic __75_D1; always_ff @(posedge aclk) begin __75_D1 <= _75; end
/*latency*/ logic __75_D2; always_ff @(posedge aclk) begin __75_D2 <= __75_D1; end
wire[15:0] _76;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _76[_g0] = value[_g0][1];
end
endgenerate
wire _77;
assign _77 = ^_76;
/*latency*/ logic __77_D1; always_ff @(posedge aclk) begin __77_D1 <= _77; end
/*latency*/ logic __77_D2; always_ff @(posedge aclk) begin __77_D2 <= __77_D1; end
wire[15:0] _78;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _78[_g0] = value[_g0][2];
end
endgenerate
wire _79;
assign _79 = ^_78;
/*latency*/ logic __79_D1; always_ff @(posedge aclk) begin __79_D1 <= _79; end
/*latency*/ logic __79_D2; always_ff @(posedge aclk) begin __79_D2 <= __79_D1; end
wire[15:0] _80;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _80[_g0] = value[_g0][3];
end
endgenerate
wire _81;
assign _81 = ^_80;
/*latency*/ logic __81_D1; always_ff @(posedge aclk) begin __81_D1 <= _81; end
/*latency*/ logic __81_D2; always_ff @(posedge aclk) begin __81_D2 <= __81_D1; end
wire[15:0] _82;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _82[_g0] = value[_g0][4];
end
endgenerate
wire _83;
assign _83 = ^_82;
/*latency*/ logic __83_D1; always_ff @(posedge aclk) begin __83_D1 <= _83; end
/*latency*/ logic __83_D2; always_ff @(posedge aclk) begin __83_D2 <= __83_D1; end
wire[15:0] _84;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _84[_g0] = value[_g0][5];
end
endgenerate
wire _85;
assign _85 = ^_84;
/*latency*/ logic __85_D1; always_ff @(posedge aclk) begin __85_D1 <= _85; end
/*latency*/ logic __85_D2; always_ff @(posedge aclk) begin __85_D2 <= __85_D1; end
wire[15:0] _86;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _86[_g0] = value[_g0][6];
end
endgenerate
wire _87;
assign _87 = ^_86;
/*latency*/ logic __87_D1; always_ff @(posedge aclk) begin __87_D1 <= _87; end
/*latency*/ logic __87_D2; always_ff @(posedge aclk) begin __87_D2 <= __87_D1; end
wire[15:0] _88;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _88[_g0] = value[_g0][7];
end
endgenerate
wire _89;
assign _89 = ^_88;
/*latency*/ logic __89_D1; always_ff @(posedge aclk) begin __89_D1 <= _89; end
/*latency*/ logic __89_D2; always_ff @(posedge aclk) begin __89_D2 <= __89_D1; end
wire[15:0] _90;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _90[_g0] = value[_g0][8];
end
endgenerate
wire _91;
assign _91 = ^_90;
/*latency*/ logic __91_D1; always_ff @(posedge aclk) begin __91_D1 <= _91; end
/*latency*/ logic __91_D2; always_ff @(posedge aclk) begin __91_D2 <= __91_D1; end
wire[15:0] _92;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _92[_g0] = value[_g0][9];
end
endgenerate
wire _93;
assign _93 = ^_92;
/*latency*/ logic __93_D1; always_ff @(posedge aclk) begin __93_D1 <= _93; end
/*latency*/ logic __93_D2; always_ff @(posedge aclk) begin __93_D2 <= __93_D1; end
wire[15:0] _94;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _94[_g0] = value[_g0][10];
end
endgenerate
wire _95;
assign _95 = ^_94;
/*latency*/ logic __95_D1; always_ff @(posedge aclk) begin __95_D1 <= _95; end
/*latency*/ logic __95_D2; always_ff @(posedge aclk) begin __95_D2 <= __95_D1; end
wire[15:0] _96;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _96[_g0] = value[_g0][11];
end
endgenerate
wire _97;
assign _97 = ^_96;
/*latency*/ logic __97_D1; always_ff @(posedge aclk) begin __97_D1 <= _97; end
/*latency*/ logic __97_D2; always_ff @(posedge aclk) begin __97_D2 <= __97_D1; end
wire[15:0] _98;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _98[_g0] = value[_g0][12];
end
endgenerate
wire _99;
assign _99 = ^_98;
/*latency*/ logic __99_D1; always_ff @(posedge aclk) begin __99_D1 <= _99; end
/*latency*/ logic __99_D2; always_ff @(posedge aclk) begin __99_D2 <= __99_D1; end
wire[15:0] _100;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _100[_g0] = value[_g0][13];
end
endgenerate
wire _101;
assign _101 = ^_100;
/*latency*/ logic __101_D1; always_ff @(posedge aclk) begin __101_D1 <= _101; end
/*latency*/ logic __101_D2; always_ff @(posedge aclk) begin __101_D2 <= __101_D1; end
wire[15:0] _102;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _102[_g0] = value[_g0][14];
end
endgenerate
wire _103;
assign _103 = ^_102;
/*latency*/ logic __103_D1; always_ff @(posedge aclk) begin __103_D1 <= _103; end
/*latency*/ logic __103_D2; always_ff @(posedge aclk) begin __103_D2 <= __103_D1; end
wire[15:0] _104;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _104[_g0] = value[_g0][15];
end
endgenerate
wire _105;
assign _105 = ^_104;
/*latency*/ logic __105_D1; always_ff @(posedge aclk) begin __105_D1 <= _105; end
/*latency*/ logic __105_D2; always_ff @(posedge aclk) begin __105_D2 <= __105_D1; end
wire[15:0] _106;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _106[_g0] = value[_g0][16];
end
endgenerate
wire _107;
assign _107 = ^_106;
/*latency*/ logic __107_D1; always_ff @(posedge aclk) begin __107_D1 <= _107; end
/*latency*/ logic __107_D2; always_ff @(posedge aclk) begin __107_D2 <= __107_D1; end
wire[15:0] _108;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _108[_g0] = value[_g0][17];
end
endgenerate
wire _109;
assign _109 = ^_108;
/*latency*/ logic __109_D1; always_ff @(posedge aclk) begin __109_D1 <= _109; end
/*latency*/ logic __109_D2; always_ff @(posedge aclk) begin __109_D2 <= __109_D1; end
wire[15:0] _110;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _110[_g0] = value[_g0][18];
end
endgenerate
wire _111;
assign _111 = ^_110;
/*latency*/ logic __111_D1; always_ff @(posedge aclk) begin __111_D1 <= _111; end
/*latency*/ logic __111_D2; always_ff @(posedge aclk) begin __111_D2 <= __111_D1; end
wire[15:0] _112;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _112[_g0] = value[_g0][19];
end
endgenerate
wire _113;
assign _113 = ^_112;
/*latency*/ logic __113_D1; always_ff @(posedge aclk) begin __113_D1 <= _113; end
/*latency*/ logic __113_D2; always_ff @(posedge aclk) begin __113_D2 <= __113_D1; end
wire[15:0] _114;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _114[_g0] = value[_g0][20];
end
endgenerate
wire _115;
assign _115 = ^_114;
/*latency*/ logic __115_D1; always_ff @(posedge aclk) begin __115_D1 <= _115; end
/*latency*/ logic __115_D2; always_ff @(posedge aclk) begin __115_D2 <= __115_D1; end
wire[15:0] _116;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _116[_g0] = value[_g0][21];
end
endgenerate
wire _117;
assign _117 = ^_116;
/*latency*/ logic __117_D1; always_ff @(posedge aclk) begin __117_D1 <= _117; end
/*latency*/ logic __117_D2; always_ff @(posedge aclk) begin __117_D2 <= __117_D1; end
wire[15:0] _118;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _118[_g0] = value[_g0][22];
end
endgenerate
wire _119;
assign _119 = ^_118;
/*latency*/ logic __119_D1; always_ff @(posedge aclk) begin __119_D1 <= _119; end
/*latency*/ logic __119_D2; always_ff @(posedge aclk) begin __119_D2 <= __119_D1; end
wire[15:0] _120;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _120[_g0] = value[_g0][23];
end
endgenerate
wire _121;
assign _121 = ^_120;
/*latency*/ logic __121_D1; always_ff @(posedge aclk) begin __121_D1 <= _121; end
/*latency*/ logic __121_D2; always_ff @(posedge aclk) begin __121_D2 <= __121_D1; end
wire[15:0] _122;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _122[_g0] = value[_g0][24];
end
endgenerate
wire _123;
assign _123 = ^_122;
/*latency*/ logic __123_D1; always_ff @(posedge aclk) begin __123_D1 <= _123; end
/*latency*/ logic __123_D2; always_ff @(posedge aclk) begin __123_D2 <= __123_D1; end
wire[15:0] _124;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _124[_g0] = value[_g0][25];
end
endgenerate
wire _125;
assign _125 = ^_124;
/*latency*/ logic __125_D1; always_ff @(posedge aclk) begin __125_D1 <= _125; end
/*latency*/ logic __125_D2; always_ff @(posedge aclk) begin __125_D2 <= __125_D1; end
wire[15:0] _126;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _126[_g0] = value[_g0][26];
end
endgenerate
wire _127;
assign _127 = ^_126;
/*latency*/ logic __127_D1; always_ff @(posedge aclk) begin __127_D1 <= _127; end
/*latency*/ logic __127_D2; always_ff @(posedge aclk) begin __127_D2 <= __127_D1; end
wire[15:0] _128;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _128[_g0] = value[_g0][27];
end
endgenerate
wire _129;
assign _129 = ^_128;
/*latency*/ logic __129_D1; always_ff @(posedge aclk) begin __129_D1 <= _129; end
/*latency*/ logic __129_D2; always_ff @(posedge aclk) begin __129_D2 <= __129_D1; end
wire[15:0] _130;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _130[_g0] = value[_g0][28];
end
endgenerate
wire _131;
assign _131 = ^_130;
/*latency*/ logic __131_D1; always_ff @(posedge aclk) begin __131_D1 <= _131; end
/*latency*/ logic __131_D2; always_ff @(posedge aclk) begin __131_D2 <= __131_D1; end
wire[15:0] _132;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _132[_g0] = value[_g0][29];
end
endgenerate
wire _133;
assign _133 = ^_132;
/*latency*/ logic __133_D1; always_ff @(posedge aclk) begin __133_D1 <= _133; end
/*latency*/ logic __133_D2; always_ff @(posedge aclk) begin __133_D2 <= __133_D1; end
wire[15:0] _134;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _134[_g0] = value[_g0][30];
end
endgenerate
wire _135;
assign _135 = ^_134;
/*latency*/ logic __135_D1; always_ff @(posedge aclk) begin __135_D1 <= _135; end
/*latency*/ logic __135_D2; always_ff @(posedge aclk) begin __135_D2 <= __135_D1; end
wire[15:0] _136;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _136[_g0] = value[_g0][31];
end
endgenerate
wire _137;
assign _137 = ^_136;
/*latency*/ logic __137_D1; always_ff @(posedge aclk) begin __137_D1 <= _137; end
/*latency*/ logic __137_D2; always_ff @(posedge aclk) begin __137_D2 <= __137_D1; end
/*mux_wire*/ logic[31:0] new_hash;
/*latency*/ logic[31:0] _new_hash_D3; always_ff @(posedge aclk) begin _new_hash_D3 <= new_hash; end
wire[31:0] _140;
assign _140 = hash ^ new_hash_contrib;
/*mux_wire*/ logic[31:0] _UIntToBits_2_value;
wire[31:0] _UIntToBits_2_bits;
/*latency*/ logic[31:0] __UIntToBits_2_bits_D1; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D1 <= _UIntToBits_2_bits; end
/*latency*/ logic[31:0] __UIntToBits_2_bits_D2; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D2 <= __UIntToBits_2_bits_D1; end
/*latency*/ logic[31:0] __UIntToBits_2_bits_D3; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D3 <= __UIntToBits_2_bits_D2; end
wire[31:0] _144;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _144[_g0] = cycles_since_reset_at_start[_g0];
end
endgenerate
wire[31:0] _145;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _145[_g0] = cycles_since_reset_at_start[32 + _g0];
end
endgenerate
wire[31:0] _146;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _146[_g0] = cycles_since_reset_bits[_g0];
end
endgenerate
wire[31:0] _147;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _147[_g0] = cycles_since_reset_bits[32 + _g0];
end
endgenerate
wire[31:0] _148[5:0];
assign _148[0] = __UIntToBits_2_bits_D3;
assign _148[1] = _new_hash_D3;
assign _148[2] = _144;
assign _148[3] = _145;
assign _148[4] = _146;
assign _148[5] = _147;
/*mux_wire*/ logic _ctrl_finish;
/*mux_wire*/ logic[31:0] _ctrl_output_regs[5:0];
wire _153;
assign _153 = !aresetn;
/*latency*/ logic __153_D1; always_ff @(posedge aclk) begin __153_D1 <= _153; end
/*latency*/ logic __153_D2; always_ff @(posedge aclk) begin __153_D2 <= __153_D1; end
localparam[31:0] _155 = 32'b00000000000000000000000000000000;
axi_ctrl_slave_NUM_INPUT_REGS_4_NUM_OUTPUT_REGS_6_ADDR_WIDTH_12_AXI_WIDTH_32 ctrl(
	.aclk(aclk),
	.aresetn(_ctrl_aresetn),
	.awaddr(_ctrl_awaddr),
	.awvalid(_ctrl_awvalid),
	.awready(_ctrl_awready),
	.wdata(_ctrl_wdata),
	.wstrb(_ctrl_wstrb),
	.wvalid(_ctrl_wvalid),
	.wready(_ctrl_wready),
	.bresp(_ctrl_bresp),
	.bvalid(_ctrl_bvalid),
	.bready(_ctrl_bready),
	.araddr(_ctrl_araddr),
	.arvalid(_ctrl_arvalid),
	.arready(_ctrl_arready),
	.rdata(_ctrl_rdata),
	.rresp(_ctrl_rresp),
	.rvalid(_ctrl_rvalid),
	.rready(_ctrl_rready),
	.input_regs(_ctrl_input_regs),
	.start(_ctrl_start),
	.finish(_ctrl_finish),
	.output_regs(_ctrl_output_regs)
);
axi_realigning_burst_reader_T_type_bool_32_16_AXI_WIDTH_512_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616 reader(
	.aclk(aclk),
	.aresetn(_reader_aresetn),
	.arvalid(_reader_arvalid),
	.arready(_reader_arready),
	.araddr(_reader_araddr),
	.arlen(_reader_arlen),
	.arsize(_reader_arsize),
	.arburst(_reader_arburst),
	.arprot(),
	.arcache(),
	.arqos(),
	.arlock(),
	.arregion(),
	.rvalid(_reader_rvalid),
	.rready(_reader_rready),
	.rdata(_reader_rdata),
	.rresp(_reader_rresp),
	.rlast(_reader_rlast),
	.max_in_flight(_reader_max_in_flight),
	.may_request_new_burst(),
	.request_new_burst(_reader_request_new_burst),
	.start_addr(_reader_start_addr),
	.count(_reader_count),
	.is_ready_to_receive_lots_of_data(_reader_is_ready_to_receive_lots_of_data),
	.value_valid(_reader_value_valid),
	.value(_reader_value),
	.last(_reader_last)
);
axi_memory_writer_tie_off_AXI_WIDTH_512 writer(
	.aclk(aclk),
	.aresetn(_writer_aresetn),
	.awvalid(_writer_awvalid),
	.awready(_writer_awready),
	.awaddr(_writer_awaddr),
	.awlen(_writer_awlen),
	.awsize(),
	.awburst(_writer_awburst),
	.awprot(),
	.awcache(_writer_awcache),
	.awqos(),
	.awlock(),
	.awregion(),
	.wvalid(_writer_wvalid),
	.wready(_writer_wready),
	.wdata(_writer_wdata),
	.wstrb(_writer_wstrb),
	.wlast(_writer_wlast),
	.bvalid(_writer_bvalid),
	.bresp(_writer_bresp),
	.bready(_writer_bready)
);
BitsToUInt_NUM_BITS_64 BitsToUInt(
	.clk(aclk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
BitsToUInt_NUM_BITS_32 BitsToUInt_2(
	.clk(aclk),
	.bits(_BitsToUInt_2_bits),
	.value(_BitsToUInt_2_value)
);
IntNarrow_FROM_I_0_TO_I_4294967296_FROM_1_TO_4294967296 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
BitsToUInt_NUM_BITS_4 BitsToUInt_3(
	.clk(aclk),
	.bits(_BitsToUInt_3_bits),
	.value(_BitsToUInt_3_value)
);
BitsToUInt_NUM_BITS_4 BitsToUInt_4(
	.clk(aclk),
	.bits(_BitsToUInt_4_bits),
	.value(_BitsToUInt_4_value)
);
BitsToUInt_NUM_BITS_11 BitsToUInt_5(
	.clk(aclk),
	.bits(_BitsToUInt_5_bits),
	.value(_BitsToUInt_5_value)
);
UIntToBits_NUM_BITS_64 UIntToBits(
	.clk(aclk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_32 UIntToBits_2(
	.clk(aclk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
always_comb begin // combinatorial _ctrl_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_aresetn = 1'bx;
	_ctrl_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_aresetn = _ctrl_aresetn;
end
always_comb begin // combinatorial s_axi_control_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_awready = 1'bx;
	s_axi_control_awready = _ctrl_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_awready = s_axi_control_awready;
end
always_comb begin // combinatorial s_axi_control_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_wready = 1'bx;
	s_axi_control_wready = _ctrl_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_wready = s_axi_control_wready;
end
always_comb begin // combinatorial s_axi_control_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bresp = 2'bxx;
	s_axi_control_bresp = _ctrl_bresp;
end
always_comb begin // combinatorial s_axi_control_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bvalid = 1'bx;
	s_axi_control_bvalid = _ctrl_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_bvalid = s_axi_control_bvalid;
end
always_comb begin // combinatorial s_axi_control_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_arready = 1'bx;
	s_axi_control_arready = _ctrl_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_arready = s_axi_control_arready;
end
always_comb begin // combinatorial s_axi_control_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	s_axi_control_rdata = _ctrl_rdata;
end
always_comb begin // combinatorial s_axi_control_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rresp = 2'bxx;
	s_axi_control_rresp = _ctrl_rresp;
end
always_comb begin // combinatorial s_axi_control_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rvalid = 1'bx;
	s_axi_control_rvalid = _ctrl_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_rvalid = s_axi_control_rvalid;
end
always_comb begin // combinatorial _ctrl_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awaddr = 12'dx;
	_ctrl_awaddr = s_axi_control_awaddr;
end
always_comb begin // combinatorial _ctrl_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awvalid = 1'bx;
	_ctrl_awvalid = s_axi_control_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_awvalid = _ctrl_awvalid;
end
always_comb begin // combinatorial _ctrl_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_ctrl_wdata = s_axi_control_wdata;
end
always_comb begin // combinatorial _ctrl_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wstrb = 4'bxxxx;
	_ctrl_wstrb = s_axi_control_wstrb;
end
always_comb begin // combinatorial _ctrl_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wvalid = 1'bx;
	_ctrl_wvalid = s_axi_control_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_wvalid = _ctrl_wvalid;
end
always_comb begin // combinatorial _ctrl_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_bready = 1'bx;
	_ctrl_bready = s_axi_control_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_bready = _ctrl_bready;
end
always_comb begin // combinatorial _ctrl_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_araddr = 12'dx;
	_ctrl_araddr = s_axi_control_araddr;
end
always_comb begin // combinatorial _ctrl_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_arvalid = 1'bx;
	_ctrl_arvalid = s_axi_control_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_arvalid = _ctrl_arvalid;
end
always_comb begin // combinatorial _ctrl_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_rready = 1'bx;
	_ctrl_rready = s_axi_control_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_rready = _ctrl_rready;
end
always_comb begin // combinatorial _reader_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_aresetn = 1'bx;
	_reader_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_aresetn = _reader_aresetn;
end
always_comb begin // combinatorial _writer_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_aresetn = 1'bx;
	_writer_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_aresetn = _writer_aresetn;
end
always_comb begin // combinatorial m_axi_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awvalid = 1'bx;
	m_axi_awvalid = _writer_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_awvalid = m_axi_awvalid;
end
always_comb begin // combinatorial m_axi_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awaddr = 64'dx;
	m_axi_awaddr = _writer_awaddr;
end
always_comb begin // combinatorial m_axi_awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awlen = 8'dx;
	m_axi_awlen = _writer_awlen;
end
always_comb begin // combinatorial m_axi_awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awburst = 2'bxx;
	m_axi_awburst = _writer_awburst;
end
always_comb begin // combinatorial m_axi_awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awcache = 4'bxxxx;
	m_axi_awcache = _writer_awcache;
end
always_comb begin // combinatorial m_axi_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wvalid = 1'bx;
	m_axi_wvalid = _writer_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wvalid = m_axi_wvalid;
end
always_comb begin // combinatorial m_axi_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wdata = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	m_axi_wdata = _writer_wdata;
end
always_comb begin // combinatorial m_axi_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wstrb = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	m_axi_wstrb = _writer_wstrb;
end
always_comb begin // combinatorial m_axi_wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wlast = 1'bx;
	m_axi_wlast = _writer_wlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wlast = m_axi_wlast;
end
always_comb begin // combinatorial m_axi_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_bready = 1'bx;
	m_axi_bready = _writer_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_bready = m_axi_bready;
end
always_comb begin // combinatorial _writer_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_awready = 1'bx;
	_writer_awready = m_axi_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_awready = _writer_awready;
end
always_comb begin // combinatorial _writer_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_wready = 1'bx;
	_writer_wready = m_axi_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_wready = _writer_wready;
end
always_comb begin // combinatorial _writer_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bvalid = 1'bx;
	_writer_bvalid = m_axi_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_bvalid = _writer_bvalid;
end
always_comb begin // combinatorial _writer_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bresp = 2'bxx;
	_writer_bresp = m_axi_bresp;
end
always_comb begin // combinatorial m_axi_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arvalid = 1'bx;
	m_axi_arvalid = _reader_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arvalid = m_axi_arvalid;
end
always_comb begin // combinatorial m_axi_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_araddr = 64'dx;
	m_axi_araddr = _reader_araddr;
end
always_comb begin // combinatorial m_axi_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlen = 8'dx;
	m_axi_arlen = _reader_arlen;
end
always_comb begin // combinatorial m_axi_arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arsize = 3'dx;
	m_axi_arsize = _reader_arsize;
end
always_comb begin // combinatorial m_axi_arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arburst = 2'bxx;
	m_axi_arburst = _reader_arburst;
end
always_comb begin // combinatorial m_axi_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_rready = 1'bx;
	m_axi_rready = _reader_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_rready = m_axi_rready;
end
always_comb begin // combinatorial _reader_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_arready = 1'bx;
	_reader_arready = m_axi_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_arready = _reader_arready;
end
always_comb begin // combinatorial _reader_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rvalid = 1'bx;
	_reader_rvalid = m_axi_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rvalid = _reader_rvalid;
end
always_comb begin // combinatorial _reader_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rdata = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_reader_rdata = m_axi_rdata;
end
always_comb begin // combinatorial _reader_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rresp = 2'bxx;
	_reader_rresp = m_axi_rresp;
end
always_comb begin // combinatorial _reader_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rlast = 1'bx;
	_reader_rlast = m_axi_rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rlast = _reader_rlast;
end
always_comb begin // combinatorial addr_a_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	addr_a_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[_v0] = _46[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[32 + _v0] = _47[_v0];
end
end
always_comb begin // combinatorial start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	start_addr = 64'dx;
	start_addr = _BitsToUInt_value;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_BitsToUInt_bits = addr_a_bits;
end
always_comb begin // combinatorial num_to_transfer
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_to_transfer = 32'dx;
	num_to_transfer = _IntNarrow_out;
end
always_comb begin // combinatorial _BitsToUInt_2_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_2_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_BitsToUInt_2_bits = _49;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 32'dx;
	_IntNarrow_in = _BitsToUInt_2_value;
end
always_comb begin // combinatorial config_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	config_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	config_bits = _50;
end
always_comb begin // combinatorial m_axi_arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arprot = 3'bxxx;
	m_axi_arprot = _51;
end
always_comb begin // combinatorial m_axi_arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arcache = 4'bxxxx;
	m_axi_arcache = _52;
end
always_comb begin // combinatorial m_axi_arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arqos = 4'dx;
	m_axi_arqos = _BitsToUInt_3_value;
end
always_comb begin // combinatorial _BitsToUInt_3_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_3_bits = 4'bxxxx;
	_BitsToUInt_3_bits = _53;
end
always_comb begin // combinatorial m_axi_arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlock = 1'bx;
	m_axi_arlock = _54;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arlock = m_axi_arlock;
end
always_comb begin // combinatorial m_axi_arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arregion = 4'dx;
	m_axi_arregion = _BitsToUInt_4_value;
end
always_comb begin // combinatorial _BitsToUInt_4_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_4_bits = 4'bxxxx;
	_BitsToUInt_4_bits = _55;
end
always_comb begin // combinatorial _BitsToUInt_5_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_5_bits = 11'bxxxxxxxxxxx;
	_BitsToUInt_5_bits = _56;
end
always_comb begin // combinatorial _reader_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_max_in_flight = 11'dx;
	_reader_max_in_flight = _BitsToUInt_5_value;
end
always_ff @(posedge aclk) begin // state cycles_since_reset
	cycles_since_reset <= _60;
	if(_153) cycles_since_reset <= 1'd0;
end
always_comb begin // combinatorial cycles_since_reset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cycles_since_reset_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	cycles_since_reset_bits = __UIntToBits_bits_D3;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 64'dx;
	_UIntToBits_value = cycles_since_reset;
end
always_ff @(posedge aclk) begin // state cycles_since_reset_at_start
	if(__ctrl_start_D3) cycles_since_reset_at_start <= cycles_since_reset_bits;
end
always_ff @(posedge aclk) begin // state running
	if(_ctrl_start) running <= 1'b1;
	if(_reader_value_valid) if(last) running <= 1'b0;
	if(_153) running <= 1'b0;
end
always_ff @(posedge aclk) begin // state num_cycles_running
	if(_ctrl_start) num_cycles_running <= 1'd0;
	if(running) num_cycles_running <= _73;
	if(_153) num_cycles_running <= 1'd0;
end
always_ff @(posedge aclk) begin // state hash
	if(__ctrl_start_D2) hash <= _67;
	if(__reader_value_valid_D2) hash <= new_hash;
	if(__153_D2) hash <= _155;
end
always_comb begin // combinatorial _reader_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_request_new_burst = 1'bx;
	_reader_request_new_burst = 1'b0;
	if(_ctrl_start) _reader_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_request_new_burst = _reader_request_new_burst;
end
always_comb begin // combinatorial _reader_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_start_addr = 64'dx;
	if(_ctrl_start) _reader_start_addr = start_addr;
end
always_comb begin // combinatorial _reader_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_count = 32'dx;
	if(_ctrl_start) _reader_count = num_to_transfer;
end
always_comb begin // combinatorial _reader_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_is_ready_to_receive_lots_of_data = 1'bx;
	_reader_is_ready_to_receive_lots_of_data = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_is_ready_to_receive_lots_of_data = _reader_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
if(_reader_value_valid) value[_v0] = _reader_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_reader_value_valid) last = _reader_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_comb begin // combinatorial new_hash_contrib
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_hash_contrib = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(__reader_value_valid_D2) new_hash_contrib[0] = __75_D2;
	if(__reader_value_valid_D2) new_hash_contrib[1] = __77_D2;
	if(__reader_value_valid_D2) new_hash_contrib[2] = __79_D2;
	if(__reader_value_valid_D2) new_hash_contrib[3] = __81_D2;
	if(__reader_value_valid_D2) new_hash_contrib[4] = __83_D2;
	if(__reader_value_valid_D2) new_hash_contrib[5] = __85_D2;
	if(__reader_value_valid_D2) new_hash_contrib[6] = __87_D2;
	if(__reader_value_valid_D2) new_hash_contrib[7] = __89_D2;
	if(__reader_value_valid_D2) new_hash_contrib[8] = __91_D2;
	if(__reader_value_valid_D2) new_hash_contrib[9] = __93_D2;
	if(__reader_value_valid_D2) new_hash_contrib[10] = __95_D2;
	if(__reader_value_valid_D2) new_hash_contrib[11] = __97_D2;
	if(__reader_value_valid_D2) new_hash_contrib[12] = __99_D2;
	if(__reader_value_valid_D2) new_hash_contrib[13] = __101_D2;
	if(__reader_value_valid_D2) new_hash_contrib[14] = __103_D2;
	if(__reader_value_valid_D2) new_hash_contrib[15] = __105_D2;
	if(__reader_value_valid_D2) new_hash_contrib[16] = __107_D2;
	if(__reader_value_valid_D2) new_hash_contrib[17] = __109_D2;
	if(__reader_value_valid_D2) new_hash_contrib[18] = __111_D2;
	if(__reader_value_valid_D2) new_hash_contrib[19] = __113_D2;
	if(__reader_value_valid_D2) new_hash_contrib[20] = __115_D2;
	if(__reader_value_valid_D2) new_hash_contrib[21] = __117_D2;
	if(__reader_value_valid_D2) new_hash_contrib[22] = __119_D2;
	if(__reader_value_valid_D2) new_hash_contrib[23] = __121_D2;
	if(__reader_value_valid_D2) new_hash_contrib[24] = __123_D2;
	if(__reader_value_valid_D2) new_hash_contrib[25] = __125_D2;
	if(__reader_value_valid_D2) new_hash_contrib[26] = __127_D2;
	if(__reader_value_valid_D2) new_hash_contrib[27] = __129_D2;
	if(__reader_value_valid_D2) new_hash_contrib[28] = __131_D2;
	if(__reader_value_valid_D2) new_hash_contrib[29] = __133_D2;
	if(__reader_value_valid_D2) new_hash_contrib[30] = __135_D2;
	if(__reader_value_valid_D2) new_hash_contrib[31] = __137_D2;
end
always_comb begin // combinatorial new_hash
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_hash = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(__reader_value_valid_D2) new_hash = _140;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 32'dx;
	if(_reader_value_valid) if(last) _UIntToBits_2_value = num_cycles_running;
end
always_comb begin // combinatorial _ctrl_finish
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_finish = 1'bx;
	_ctrl_finish = 1'b0;
	if(__reader_value_valid_D3) if(_last_D3) _ctrl_finish = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_finish = _ctrl_finish;
end
always_comb begin // combinatorial _ctrl_output_regs
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_output_regs = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
if(__reader_value_valid_D3) if(_last_D3) _ctrl_output_regs[_v0] = _148[_v0];
end
end
endmodule

// axi_memory_writer_tie_off #(AXI_WIDTH: 512)
module axi_memory_writer_tie_off_AXI_WIDTH_512(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic awvalid,
	input wire awready,
	output /*mux_wire*/ logic[63:0] awaddr,
	output /*mux_wire*/ logic[7:0] awlen,
	output /*mux_wire*/ logic[2:0] awsize,
	output /*mux_wire*/ logic[1:0] awburst,
	output /*mux_wire*/ logic[2:0] awprot,
	output /*mux_wire*/ logic[3:0] awcache,
	output /*mux_wire*/ logic[3:0] awqos,
	output /*mux_wire*/ logic awlock,
	output /*mux_wire*/ logic[3:0] awregion,
	output /*mux_wire*/ logic wvalid,
	input wire wready,
	output /*mux_wire*/ logic[511:0] wdata,
	output /*mux_wire*/ logic[63:0] wstrb,
	output /*mux_wire*/ logic wlast,
	input wire bvalid,
	input wire[1:0] bresp,
	output /*mux_wire*/ logic bready
);

/*mux_wire*/ logic _aresetn;
localparam[1:0] _4 = 2'b00;
localparam[2:0] _5 = 3'b000;
localparam[3:0] _6 = 4'b0000;
/*mux_wire*/ logic _Repeat_v;
wire[511:0] _Repeat_result;
/*mux_wire*/ logic _Repeat_2_v;
wire[63:0] _Repeat_2_result;
/*mux_wire*/ logic _awready;
/*mux_wire*/ logic _wready;
/*mux_wire*/ logic _bvalid;
/*mux_wire*/ logic[1:0] _bresp;
Repeat_T_type_bool_SIZE_512 Repeat(
	.clk(aclk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
Repeat_T_type_bool_SIZE_64 Repeat_2(
	.clk(aclk),
	.v(_Repeat_2_v),
	.result(_Repeat_2_result)
);
always_comb begin // combinatorial _aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_aresetn = 1'bx;
	_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_aresetn = _aresetn;
end
always_comb begin // combinatorial awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awvalid = 1'bx;
	awvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awvalid = awvalid;
end
always_comb begin // combinatorial awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awaddr = 64'dx;
	awaddr = 1'd0;
end
always_comb begin // combinatorial awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlen = 8'dx;
	awlen = 1'd0;
end
always_comb begin // combinatorial awsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awsize = 3'dx;
	awsize = 3'd6;
end
always_comb begin // combinatorial awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awburst = 2'bxx;
	awburst = _4;
end
always_comb begin // combinatorial awprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awprot = 3'bxxx;
	awprot = _5;
end
always_comb begin // combinatorial awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awcache = 4'bxxxx;
	awcache = _6;
end
always_comb begin // combinatorial awqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awqos = 4'dx;
	awqos = 1'd0;
end
always_comb begin // combinatorial awlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlock = 1'bx;
	awlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awlock = awlock;
end
always_comb begin // combinatorial awregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awregion = 4'dx;
	awregion = 1'd0;
end
always_comb begin // combinatorial wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wvalid = 1'bx;
	wvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wvalid = wvalid;
end
always_comb begin // combinatorial wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wdata = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	wdata = _Repeat_result;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	_Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
always_comb begin // combinatorial wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wstrb = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	wstrb = _Repeat_2_result;
end
always_comb begin // combinatorial _Repeat_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_2_v = 1'bx;
	_Repeat_2_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_2_v = _Repeat_2_v;
end
always_comb begin // combinatorial wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wlast = 1'bx;
	wlast = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wlast = wlast;
end
always_comb begin // combinatorial bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	bready = 1'bx;
	bready = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	bready = bready;
end
always_comb begin // combinatorial _awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_awready = 1'bx;
	_awready = awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_awready = _awready;
end
always_comb begin // combinatorial _wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_wready = 1'bx;
	_wready = wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_wready = _wready;
end
always_comb begin // combinatorial _bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_bvalid = 1'bx;
	_bvalid = bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_bvalid = _bvalid;
end
always_comb begin // combinatorial _bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_bresp = 2'bxx;
	_bresp = bresp;
end
endmodule

// Repeat #(T: type bool #(), SIZE: 512)
module Repeat_T_type_bool_SIZE_512(
	input clk,
	input wire v,
	output /*mux_wire*/ logic[511:0] result
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
	result[4] = v;
	result[5] = v;
	result[6] = v;
	result[7] = v;
	result[8] = v;
	result[9] = v;
	result[10] = v;
	result[11] = v;
	result[12] = v;
	result[13] = v;
	result[14] = v;
	result[15] = v;
	result[16] = v;
	result[17] = v;
	result[18] = v;
	result[19] = v;
	result[20] = v;
	result[21] = v;
	result[22] = v;
	result[23] = v;
	result[24] = v;
	result[25] = v;
	result[26] = v;
	result[27] = v;
	result[28] = v;
	result[29] = v;
	result[30] = v;
	result[31] = v;
	result[32] = v;
	result[33] = v;
	result[34] = v;
	result[35] = v;
	result[36] = v;
	result[37] = v;
	result[38] = v;
	result[39] = v;
	result[40] = v;
	result[41] = v;
	result[42] = v;
	result[43] = v;
	result[44] = v;
	result[45] = v;
	result[46] = v;
	result[47] = v;
	result[48] = v;
	result[49] = v;
	result[50] = v;
	result[51] = v;
	result[52] = v;
	result[53] = v;
	result[54] = v;
	result[55] = v;
	result[56] = v;
	result[57] = v;
	result[58] = v;
	result[59] = v;
	result[60] = v;
	result[61] = v;
	result[62] = v;
	result[63] = v;
	result[64] = v;
	result[65] = v;
	result[66] = v;
	result[67] = v;
	result[68] = v;
	result[69] = v;
	result[70] = v;
	result[71] = v;
	result[72] = v;
	result[73] = v;
	result[74] = v;
	result[75] = v;
	result[76] = v;
	result[77] = v;
	result[78] = v;
	result[79] = v;
	result[80] = v;
	result[81] = v;
	result[82] = v;
	result[83] = v;
	result[84] = v;
	result[85] = v;
	result[86] = v;
	result[87] = v;
	result[88] = v;
	result[89] = v;
	result[90] = v;
	result[91] = v;
	result[92] = v;
	result[93] = v;
	result[94] = v;
	result[95] = v;
	result[96] = v;
	result[97] = v;
	result[98] = v;
	result[99] = v;
	result[100] = v;
	result[101] = v;
	result[102] = v;
	result[103] = v;
	result[104] = v;
	result[105] = v;
	result[106] = v;
	result[107] = v;
	result[108] = v;
	result[109] = v;
	result[110] = v;
	result[111] = v;
	result[112] = v;
	result[113] = v;
	result[114] = v;
	result[115] = v;
	result[116] = v;
	result[117] = v;
	result[118] = v;
	result[119] = v;
	result[120] = v;
	result[121] = v;
	result[122] = v;
	result[123] = v;
	result[124] = v;
	result[125] = v;
	result[126] = v;
	result[127] = v;
	result[128] = v;
	result[129] = v;
	result[130] = v;
	result[131] = v;
	result[132] = v;
	result[133] = v;
	result[134] = v;
	result[135] = v;
	result[136] = v;
	result[137] = v;
	result[138] = v;
	result[139] = v;
	result[140] = v;
	result[141] = v;
	result[142] = v;
	result[143] = v;
	result[144] = v;
	result[145] = v;
	result[146] = v;
	result[147] = v;
	result[148] = v;
	result[149] = v;
	result[150] = v;
	result[151] = v;
	result[152] = v;
	result[153] = v;
	result[154] = v;
	result[155] = v;
	result[156] = v;
	result[157] = v;
	result[158] = v;
	result[159] = v;
	result[160] = v;
	result[161] = v;
	result[162] = v;
	result[163] = v;
	result[164] = v;
	result[165] = v;
	result[166] = v;
	result[167] = v;
	result[168] = v;
	result[169] = v;
	result[170] = v;
	result[171] = v;
	result[172] = v;
	result[173] = v;
	result[174] = v;
	result[175] = v;
	result[176] = v;
	result[177] = v;
	result[178] = v;
	result[179] = v;
	result[180] = v;
	result[181] = v;
	result[182] = v;
	result[183] = v;
	result[184] = v;
	result[185] = v;
	result[186] = v;
	result[187] = v;
	result[188] = v;
	result[189] = v;
	result[190] = v;
	result[191] = v;
	result[192] = v;
	result[193] = v;
	result[194] = v;
	result[195] = v;
	result[196] = v;
	result[197] = v;
	result[198] = v;
	result[199] = v;
	result[200] = v;
	result[201] = v;
	result[202] = v;
	result[203] = v;
	result[204] = v;
	result[205] = v;
	result[206] = v;
	result[207] = v;
	result[208] = v;
	result[209] = v;
	result[210] = v;
	result[211] = v;
	result[212] = v;
	result[213] = v;
	result[214] = v;
	result[215] = v;
	result[216] = v;
	result[217] = v;
	result[218] = v;
	result[219] = v;
	result[220] = v;
	result[221] = v;
	result[222] = v;
	result[223] = v;
	result[224] = v;
	result[225] = v;
	result[226] = v;
	result[227] = v;
	result[228] = v;
	result[229] = v;
	result[230] = v;
	result[231] = v;
	result[232] = v;
	result[233] = v;
	result[234] = v;
	result[235] = v;
	result[236] = v;
	result[237] = v;
	result[238] = v;
	result[239] = v;
	result[240] = v;
	result[241] = v;
	result[242] = v;
	result[243] = v;
	result[244] = v;
	result[245] = v;
	result[246] = v;
	result[247] = v;
	result[248] = v;
	result[249] = v;
	result[250] = v;
	result[251] = v;
	result[252] = v;
	result[253] = v;
	result[254] = v;
	result[255] = v;
	result[256] = v;
	result[257] = v;
	result[258] = v;
	result[259] = v;
	result[260] = v;
	result[261] = v;
	result[262] = v;
	result[263] = v;
	result[264] = v;
	result[265] = v;
	result[266] = v;
	result[267] = v;
	result[268] = v;
	result[269] = v;
	result[270] = v;
	result[271] = v;
	result[272] = v;
	result[273] = v;
	result[274] = v;
	result[275] = v;
	result[276] = v;
	result[277] = v;
	result[278] = v;
	result[279] = v;
	result[280] = v;
	result[281] = v;
	result[282] = v;
	result[283] = v;
	result[284] = v;
	result[285] = v;
	result[286] = v;
	result[287] = v;
	result[288] = v;
	result[289] = v;
	result[290] = v;
	result[291] = v;
	result[292] = v;
	result[293] = v;
	result[294] = v;
	result[295] = v;
	result[296] = v;
	result[297] = v;
	result[298] = v;
	result[299] = v;
	result[300] = v;
	result[301] = v;
	result[302] = v;
	result[303] = v;
	result[304] = v;
	result[305] = v;
	result[306] = v;
	result[307] = v;
	result[308] = v;
	result[309] = v;
	result[310] = v;
	result[311] = v;
	result[312] = v;
	result[313] = v;
	result[314] = v;
	result[315] = v;
	result[316] = v;
	result[317] = v;
	result[318] = v;
	result[319] = v;
	result[320] = v;
	result[321] = v;
	result[322] = v;
	result[323] = v;
	result[324] = v;
	result[325] = v;
	result[326] = v;
	result[327] = v;
	result[328] = v;
	result[329] = v;
	result[330] = v;
	result[331] = v;
	result[332] = v;
	result[333] = v;
	result[334] = v;
	result[335] = v;
	result[336] = v;
	result[337] = v;
	result[338] = v;
	result[339] = v;
	result[340] = v;
	result[341] = v;
	result[342] = v;
	result[343] = v;
	result[344] = v;
	result[345] = v;
	result[346] = v;
	result[347] = v;
	result[348] = v;
	result[349] = v;
	result[350] = v;
	result[351] = v;
	result[352] = v;
	result[353] = v;
	result[354] = v;
	result[355] = v;
	result[356] = v;
	result[357] = v;
	result[358] = v;
	result[359] = v;
	result[360] = v;
	result[361] = v;
	result[362] = v;
	result[363] = v;
	result[364] = v;
	result[365] = v;
	result[366] = v;
	result[367] = v;
	result[368] = v;
	result[369] = v;
	result[370] = v;
	result[371] = v;
	result[372] = v;
	result[373] = v;
	result[374] = v;
	result[375] = v;
	result[376] = v;
	result[377] = v;
	result[378] = v;
	result[379] = v;
	result[380] = v;
	result[381] = v;
	result[382] = v;
	result[383] = v;
	result[384] = v;
	result[385] = v;
	result[386] = v;
	result[387] = v;
	result[388] = v;
	result[389] = v;
	result[390] = v;
	result[391] = v;
	result[392] = v;
	result[393] = v;
	result[394] = v;
	result[395] = v;
	result[396] = v;
	result[397] = v;
	result[398] = v;
	result[399] = v;
	result[400] = v;
	result[401] = v;
	result[402] = v;
	result[403] = v;
	result[404] = v;
	result[405] = v;
	result[406] = v;
	result[407] = v;
	result[408] = v;
	result[409] = v;
	result[410] = v;
	result[411] = v;
	result[412] = v;
	result[413] = v;
	result[414] = v;
	result[415] = v;
	result[416] = v;
	result[417] = v;
	result[418] = v;
	result[419] = v;
	result[420] = v;
	result[421] = v;
	result[422] = v;
	result[423] = v;
	result[424] = v;
	result[425] = v;
	result[426] = v;
	result[427] = v;
	result[428] = v;
	result[429] = v;
	result[430] = v;
	result[431] = v;
	result[432] = v;
	result[433] = v;
	result[434] = v;
	result[435] = v;
	result[436] = v;
	result[437] = v;
	result[438] = v;
	result[439] = v;
	result[440] = v;
	result[441] = v;
	result[442] = v;
	result[443] = v;
	result[444] = v;
	result[445] = v;
	result[446] = v;
	result[447] = v;
	result[448] = v;
	result[449] = v;
	result[450] = v;
	result[451] = v;
	result[452] = v;
	result[453] = v;
	result[454] = v;
	result[455] = v;
	result[456] = v;
	result[457] = v;
	result[458] = v;
	result[459] = v;
	result[460] = v;
	result[461] = v;
	result[462] = v;
	result[463] = v;
	result[464] = v;
	result[465] = v;
	result[466] = v;
	result[467] = v;
	result[468] = v;
	result[469] = v;
	result[470] = v;
	result[471] = v;
	result[472] = v;
	result[473] = v;
	result[474] = v;
	result[475] = v;
	result[476] = v;
	result[477] = v;
	result[478] = v;
	result[479] = v;
	result[480] = v;
	result[481] = v;
	result[482] = v;
	result[483] = v;
	result[484] = v;
	result[485] = v;
	result[486] = v;
	result[487] = v;
	result[488] = v;
	result[489] = v;
	result[490] = v;
	result[491] = v;
	result[492] = v;
	result[493] = v;
	result[494] = v;
	result[495] = v;
	result[496] = v;
	result[497] = v;
	result[498] = v;
	result[499] = v;
	result[500] = v;
	result[501] = v;
	result[502] = v;
	result[503] = v;
	result[504] = v;
	result[505] = v;
	result[506] = v;
	result[507] = v;
	result[508] = v;
	result[509] = v;
	result[510] = v;
	result[511] = v;
end
endmodule

// axi_realigning_burst_reader #(T: type bool #()[32][16], AXI_WIDTH: 512, ADDR_ALIGN: 4, COUNT_TO: 4294967296, ATO: 18446744073709551616)
module axi_realigning_burst_reader_T_type_bool_32_16_AXI_WIDTH_512_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic arvalid,
	input wire arready,
	output /*mux_wire*/ logic[63:0] araddr,
	output /*mux_wire*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[511:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[31:0] count,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic value_valid,
	output /*mux_wire*/ logic[31:0] value[15:0],
	output /*mux_wire*/ logic last
);

/*mux_wire*/ logic _parent_aresetn;
wire _parent_arvalid;
wire[63:0] _parent_araddr;
wire[7:0] _parent_arlen;
wire[2:0] _parent_arsize;
wire[1:0] _parent_arburst;
wire[2:0] _parent_arprot;
wire[3:0] _parent_arcache;
wire[3:0] _parent_arqos;
wire _parent_arlock;
wire[3:0] _parent_arregion;
wire _parent_rready;
/*mux_wire*/ logic _parent_arready;
/*mux_wire*/ logic _parent_rvalid;
/*mux_wire*/ logic[511:0] _parent_rdata;
/*mux_wire*/ logic[1:0] _parent_rresp;
/*mux_wire*/ logic _parent_rlast;
/*mux_wire*/ logic[10:0] _parent_max_in_flight;
wire _parent_may_request_new_burst;
wire[35:0] _22;
assign _22 = count * 5'd16;
/*mux_wire*/ logic _parent_request_new_burst;
/*mux_wire*/ logic[63:0] _parent_start_addr;
/*mux_wire*/ logic[35:0] _parent_count;
/*mux_wire*/ logic _parent_is_ready_to_receive_lots_of_data;
/*state*/ logic[31:0] stored_elements[14:0];
/*state*/ logic[3:0] cur_element_store_align;
wire _parent_element_packet_valid;
wire[31:0] _parent_elements[15:0];
wire[3:0] _parent_chunk_offset;
wire[4:0] _parent_chunk_length;
wire _parent_last;
/*mux_wire*/ logic[31:0] elements[15:0];
/*mux_wire*/ logic[3:0] chunk_offset;
/*mux_wire*/ logic[4:0] chunk_length;
/*mux_wire*/ logic last_2;
/*mux_wire*/ logic[31:0] elements_extended[15:0];
/*mux_wire*/ logic[31:0] rotated_elements[15:0];
wire signed[4:0] _31;
assign _31 = cur_element_store_align - chunk_offset;
wire[3:0] _32;
assign _32 = _31; // == mod 16 (target is 4 bits wide)
/*mux_wire*/ logic[31:0] _RotateRight_data[15:0];
/*mux_wire*/ logic[3:0] _RotateRight_offset;
wire[31:0] _RotateRight_rotated_data[15:0];
/*mux_wire*/ logic[15:0] rotated_strobe;
/*mux_wire*/ logic[3:0] _MakeStrobe_chunk_offset;
/*mux_wire*/ logic[4:0] _MakeStrobe_chunk_length;
wire[15:0] _MakeStrobe_strobe;
/*mux_wire*/ logic[4:0] end_of_element;
wire[4:0] _37;
assign _37 = cur_element_store_align + chunk_length;
wire _39;
assign _39 = end_of_element >= 5'd16;
/*mux_wire*/ logic[511:0] resulting_value_bits;
wire _41;
assign _41 = cur_element_store_align > 1'd0;
wire[31:0] _42 = stored_elements[0];
wire[31:0] _43 = rotated_elements[0];
wire _45;
assign _45 = cur_element_store_align > 1'd1;
wire[31:0] _46 = stored_elements[1];
wire[31:0] _47 = rotated_elements[1];
wire _49;
assign _49 = cur_element_store_align > 2'd2;
wire[31:0] _50 = stored_elements[2];
wire[31:0] _51 = rotated_elements[2];
wire _53;
assign _53 = cur_element_store_align > 2'd3;
wire[31:0] _54 = stored_elements[3];
wire[31:0] _55 = rotated_elements[3];
wire _57;
assign _57 = cur_element_store_align > 3'd4;
wire[31:0] _58 = stored_elements[4];
wire[31:0] _59 = rotated_elements[4];
wire _61;
assign _61 = cur_element_store_align > 3'd5;
wire[31:0] _62 = stored_elements[5];
wire[31:0] _63 = rotated_elements[5];
wire _65;
assign _65 = cur_element_store_align > 3'd6;
wire[31:0] _66 = stored_elements[6];
wire[31:0] _67 = rotated_elements[6];
wire _69;
assign _69 = cur_element_store_align > 3'd7;
wire[31:0] _70 = stored_elements[7];
wire[31:0] _71 = rotated_elements[7];
wire _73;
assign _73 = cur_element_store_align > 4'd8;
wire[31:0] _74 = stored_elements[8];
wire[31:0] _75 = rotated_elements[8];
wire _77;
assign _77 = cur_element_store_align > 4'd9;
wire[31:0] _78 = stored_elements[9];
wire[31:0] _79 = rotated_elements[9];
wire _81;
assign _81 = cur_element_store_align > 4'd10;
wire[31:0] _82 = stored_elements[10];
wire[31:0] _83 = rotated_elements[10];
wire _85;
assign _85 = cur_element_store_align > 4'd11;
wire[31:0] _86 = stored_elements[11];
wire[31:0] _87 = rotated_elements[11];
wire _89;
assign _89 = cur_element_store_align > 4'd12;
wire[31:0] _90 = stored_elements[12];
wire[31:0] _91 = rotated_elements[12];
wire _93;
assign _93 = cur_element_store_align > 4'd13;
wire[31:0] _94 = stored_elements[13];
wire[31:0] _95 = rotated_elements[13];
wire _97;
assign _97 = cur_element_store_align > 4'd14;
wire[31:0] _98 = stored_elements[14];
wire[31:0] _99 = rotated_elements[14];
wire[31:0] _100 = rotated_elements[15];
/*mux_wire*/ logic[511:0] _FromBits_bits;
wire[31:0] _FromBits_value[15:0];
wire[3:0] _105;
assign _105 = end_of_element; // == mod 16 (target is 4 bits wide)
wire _106 = rotated_strobe[0];
wire[31:0] _107 = rotated_elements[0];
wire _108 = rotated_strobe[1];
wire[31:0] _109 = rotated_elements[1];
wire _110 = rotated_strobe[2];
wire[31:0] _111 = rotated_elements[2];
wire _112 = rotated_strobe[3];
wire[31:0] _113 = rotated_elements[3];
wire _114 = rotated_strobe[4];
wire[31:0] _115 = rotated_elements[4];
wire _116 = rotated_strobe[5];
wire[31:0] _117 = rotated_elements[5];
wire _118 = rotated_strobe[6];
wire[31:0] _119 = rotated_elements[6];
wire _120 = rotated_strobe[7];
wire[31:0] _121 = rotated_elements[7];
wire _122 = rotated_strobe[8];
wire[31:0] _123 = rotated_elements[8];
wire _124 = rotated_strobe[9];
wire[31:0] _125 = rotated_elements[9];
wire _126 = rotated_strobe[10];
wire[31:0] _127 = rotated_elements[10];
wire _128 = rotated_strobe[11];
wire[31:0] _129 = rotated_elements[11];
wire _130 = rotated_strobe[12];
wire[31:0] _131 = rotated_elements[12];
wire _132 = rotated_strobe[13];
wire[31:0] _133 = rotated_elements[13];
wire _134 = rotated_strobe[14];
wire[31:0] _135 = rotated_elements[14];
wire _137;
assign _137 = !aresetn;
axi_array_burst_reader_AXI_WIDTH_512_ADDR_ALIGN_4_COUNT_TO_68719476736_ATO_18446744073709551616 parent(
	.aclk(aclk),
	.aresetn(_parent_aresetn),
	.arvalid(_parent_arvalid),
	.arready(_parent_arready),
	.araddr(_parent_araddr),
	.arlen(_parent_arlen),
	.arsize(_parent_arsize),
	.arburst(_parent_arburst),
	.arprot(_parent_arprot),
	.arcache(_parent_arcache),
	.arqos(_parent_arqos),
	.arlock(_parent_arlock),
	.arregion(_parent_arregion),
	.rvalid(_parent_rvalid),
	.rready(_parent_rready),
	.rdata(_parent_rdata),
	.rresp(_parent_rresp),
	.rlast(_parent_rlast),
	.is_ready_to_receive_lots_of_data(_parent_is_ready_to_receive_lots_of_data),
	.element_packet_valid(_parent_element_packet_valid),
	.elements(_parent_elements),
	.chunk_offset(_parent_chunk_offset),
	.chunk_length(_parent_chunk_length),
	.last(_parent_last),
	.max_in_flight(_parent_max_in_flight),
	.may_request_new_burst(_parent_may_request_new_burst),
	.request_new_burst(_parent_request_new_burst),
	.start_addr(_parent_start_addr),
	.count(_parent_count)
);
RotateRight_T_type_bool_32_ARRAY_LEN_16 RotateRight(
	.clk(aclk),
	.data(_RotateRight_data),
	.offset(_RotateRight_offset),
	.rotated_data(_RotateRight_rotated_data)
);
MakeStrobe_STROBE_WIDTH_16 MakeStrobe(
	.clk(aclk),
	.chunk_offset(_MakeStrobe_chunk_offset),
	.chunk_length(_MakeStrobe_chunk_length),
	.strobe(_MakeStrobe_strobe)
);
FromBits_T_type_bool_32_16 FromBits(
	.clk(aclk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial _parent_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_aresetn = 1'bx;
	_parent_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_aresetn = _parent_aresetn;
end
always_comb begin // combinatorial arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arvalid = 1'bx;
	arvalid = _parent_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arvalid = arvalid;
end
always_comb begin // combinatorial araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	araddr = 64'dx;
	araddr = _parent_araddr;
end
always_comb begin // combinatorial arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlen = 8'dx;
	arlen = _parent_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = _parent_arsize;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _parent_arburst;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _parent_arprot;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _parent_arcache;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = _parent_arqos;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = _parent_arlock;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = _parent_arregion;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = _parent_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _parent_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_arready = 1'bx;
	_parent_arready = arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_arready = _parent_arready;
end
always_comb begin // combinatorial _parent_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rvalid = 1'bx;
	_parent_rvalid = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rvalid = _parent_rvalid;
end
always_comb begin // combinatorial _parent_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rdata = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_parent_rdata = rdata;
end
always_comb begin // combinatorial _parent_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rresp = 2'bxx;
	_parent_rresp = rresp;
end
always_comb begin // combinatorial _parent_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rlast = 1'bx;
	_parent_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rlast = _parent_rlast;
end
always_comb begin // combinatorial _parent_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_max_in_flight = 11'dx;
	_parent_max_in_flight = max_in_flight;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _parent_may_request_new_burst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial _parent_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_request_new_burst = 1'bx;
	_parent_request_new_burst = 1'b0;
	if(request_new_burst) _parent_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_request_new_burst = _parent_request_new_burst;
end
always_comb begin // combinatorial _parent_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_start_addr = 64'dx;
	if(request_new_burst) _parent_start_addr = start_addr;
end
always_comb begin // combinatorial _parent_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_count = 36'dx;
	if(request_new_burst) _parent_count = _22;
end
always_comb begin // combinatorial _parent_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_is_ready_to_receive_lots_of_data = 1'bx;
	_parent_is_ready_to_receive_lots_of_data = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_is_ready_to_receive_lots_of_data = _parent_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value_valid = 1'bx;
	value_valid = 1'b0;
	if(_parent_element_packet_valid) if(_39) value_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	value_valid = value_valid;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) value[_v0] = _FromBits_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_parent_element_packet_valid) if(_39) last = last_2;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state stored_elements
	if(_parent_element_packet_valid) if(_106) stored_elements[0] <= _107;
	if(_parent_element_packet_valid) if(_108) stored_elements[1] <= _109;
	if(_parent_element_packet_valid) if(_110) stored_elements[2] <= _111;
	if(_parent_element_packet_valid) if(_112) stored_elements[3] <= _113;
	if(_parent_element_packet_valid) if(_114) stored_elements[4] <= _115;
	if(_parent_element_packet_valid) if(_116) stored_elements[5] <= _117;
	if(_parent_element_packet_valid) if(_118) stored_elements[6] <= _119;
	if(_parent_element_packet_valid) if(_120) stored_elements[7] <= _121;
	if(_parent_element_packet_valid) if(_122) stored_elements[8] <= _123;
	if(_parent_element_packet_valid) if(_124) stored_elements[9] <= _125;
	if(_parent_element_packet_valid) if(_126) stored_elements[10] <= _127;
	if(_parent_element_packet_valid) if(_128) stored_elements[11] <= _129;
	if(_parent_element_packet_valid) if(_130) stored_elements[12] <= _131;
	if(_parent_element_packet_valid) if(_132) stored_elements[13] <= _133;
	if(_parent_element_packet_valid) if(_134) stored_elements[14] <= _135;
end
always_ff @(posedge aclk) begin // state cur_element_store_align
	if(_parent_element_packet_valid) cur_element_store_align <= _105;
	if(_137) cur_element_store_align <= 1'd0;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements[_v0] = _parent_elements[_v0];
end
end
always_comb begin // combinatorial chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_offset = 4'dx;
	if(_parent_element_packet_valid) chunk_offset = _parent_chunk_offset;
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 5'dx;
	if(_parent_element_packet_valid) chunk_length = _parent_chunk_length;
end
always_comb begin // combinatorial last_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last_2 = 1'bx;
	if(_parent_element_packet_valid) last_2 = _parent_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last_2 = last_2;
end
always_comb begin // combinatorial elements_extended
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_extended = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements_extended[_v0] = elements[_v0];
end
end
always_comb begin // combinatorial rotated_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) rotated_elements[_v0] = _RotateRight_rotated_data[_v0];
end
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) _RotateRight_data[_v0] = elements_extended[_v0];
end
end
always_comb begin // combinatorial _RotateRight_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_offset = 4'dx;
	if(_parent_element_packet_valid) _RotateRight_offset = _32;
end
always_comb begin // combinatorial rotated_strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_strobe = 16'bxxxxxxxxxxxxxxxx;
	if(_parent_element_packet_valid) rotated_strobe = _MakeStrobe_strobe;
end
always_comb begin // combinatorial _MakeStrobe_chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_offset = 4'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_offset = cur_element_store_align;
end
always_comb begin // combinatorial _MakeStrobe_chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_length = 5'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_length = chunk_length;
end
always_comb begin // combinatorial end_of_element
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	end_of_element = 5'dx;
	if(_parent_element_packet_valid) end_of_element = _37;
end
always_comb begin // combinatorial resulting_value_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	resulting_value_bits = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_41) resulting_value_bits[_v0] = _42[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_41) resulting_value_bits[_v0] = _43[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_45) resulting_value_bits[32 + _v0] = _46[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_45) resulting_value_bits[32 + _v0] = _47[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_49) resulting_value_bits[64 + _v0] = _50[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_49) resulting_value_bits[64 + _v0] = _51[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_53) resulting_value_bits[96 + _v0] = _54[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_53) resulting_value_bits[96 + _v0] = _55[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_57) resulting_value_bits[128 + _v0] = _58[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_57) resulting_value_bits[128 + _v0] = _59[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_61) resulting_value_bits[160 + _v0] = _62[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_61) resulting_value_bits[160 + _v0] = _63[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_65) resulting_value_bits[192 + _v0] = _66[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_65) resulting_value_bits[192 + _v0] = _67[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_69) resulting_value_bits[224 + _v0] = _70[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_69) resulting_value_bits[224 + _v0] = _71[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_73) resulting_value_bits[256 + _v0] = _74[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_73) resulting_value_bits[256 + _v0] = _75[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_77) resulting_value_bits[288 + _v0] = _78[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_77) resulting_value_bits[288 + _v0] = _79[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_81) resulting_value_bits[320 + _v0] = _82[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_81) resulting_value_bits[320 + _v0] = _83[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_85) resulting_value_bits[352 + _v0] = _86[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_85) resulting_value_bits[352 + _v0] = _87[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_89) resulting_value_bits[384 + _v0] = _90[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_89) resulting_value_bits[384 + _v0] = _91[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_93) resulting_value_bits[416 + _v0] = _94[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_93) resulting_value_bits[416 + _v0] = _95[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_97) resulting_value_bits[448 + _v0] = _98[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_97) resulting_value_bits[448 + _v0] = _99[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) resulting_value_bits[480 + _v0] = _100[_v0];
end
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_parent_element_packet_valid) if(_39) _FromBits_bits = resulting_value_bits;
end
endmodule

// MakeStrobe #(STROBE_WIDTH: 16)
module MakeStrobe_STROBE_WIDTH_16(
	input clk,
	input wire[3:0] chunk_offset,
	input wire[4:0] chunk_length,
	output /*mux_wire*/ logic[15:0] strobe
);

/*mux_wire*/ logic[15:0] chunk_bits;
wire _2;
assign _2 = chunk_length > 1'd0;
wire _4;
assign _4 = chunk_length > 1'd1;
wire _6;
assign _6 = chunk_length > 2'd2;
wire _8;
assign _8 = chunk_length > 2'd3;
wire _10;
assign _10 = chunk_length > 3'd4;
wire _12;
assign _12 = chunk_length > 3'd5;
wire _14;
assign _14 = chunk_length > 3'd6;
wire _16;
assign _16 = chunk_length > 3'd7;
wire _18;
assign _18 = chunk_length > 4'd8;
wire _20;
assign _20 = chunk_length > 4'd9;
wire _22;
assign _22 = chunk_length > 4'd10;
wire _24;
assign _24 = chunk_length > 4'd11;
wire _26;
assign _26 = chunk_length > 4'd12;
wire _28;
assign _28 = chunk_length > 4'd13;
wire _30;
assign _30 = chunk_length > 4'd14;
wire _32;
assign _32 = chunk_length > 4'd15;
/*mux_wire*/ logic[15:0] _RotateRight_data;
/*mux_wire*/ logic[3:0] _RotateRight_offset;
wire[15:0] _RotateRight_rotated_data;
RotateRight_T_type_bool_ARRAY_LEN_16 RotateRight(
	.clk(clk),
	.data(_RotateRight_data),
	.offset(_RotateRight_offset),
	.rotated_data(_RotateRight_rotated_data)
);
always_comb begin // combinatorial strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	strobe = 16'bxxxxxxxxxxxxxxxx;
	strobe = _RotateRight_rotated_data;
end
always_comb begin // combinatorial chunk_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_bits = 16'bxxxxxxxxxxxxxxxx;
	if(_2) chunk_bits[0] = 1'b1;
	if(!_2) chunk_bits[0] = 1'b0;
	if(_4) chunk_bits[1] = 1'b1;
	if(!_4) chunk_bits[1] = 1'b0;
	if(_6) chunk_bits[2] = 1'b1;
	if(!_6) chunk_bits[2] = 1'b0;
	if(_8) chunk_bits[3] = 1'b1;
	if(!_8) chunk_bits[3] = 1'b0;
	if(_10) chunk_bits[4] = 1'b1;
	if(!_10) chunk_bits[4] = 1'b0;
	if(_12) chunk_bits[5] = 1'b1;
	if(!_12) chunk_bits[5] = 1'b0;
	if(_14) chunk_bits[6] = 1'b1;
	if(!_14) chunk_bits[6] = 1'b0;
	if(_16) chunk_bits[7] = 1'b1;
	if(!_16) chunk_bits[7] = 1'b0;
	if(_18) chunk_bits[8] = 1'b1;
	if(!_18) chunk_bits[8] = 1'b0;
	if(_20) chunk_bits[9] = 1'b1;
	if(!_20) chunk_bits[9] = 1'b0;
	if(_22) chunk_bits[10] = 1'b1;
	if(!_22) chunk_bits[10] = 1'b0;
	if(_24) chunk_bits[11] = 1'b1;
	if(!_24) chunk_bits[11] = 1'b0;
	if(_26) chunk_bits[12] = 1'b1;
	if(!_26) chunk_bits[12] = 1'b0;
	if(_28) chunk_bits[13] = 1'b1;
	if(!_28) chunk_bits[13] = 1'b0;
	if(_30) chunk_bits[14] = 1'b1;
	if(!_30) chunk_bits[14] = 1'b0;
	if(_32) chunk_bits[15] = 1'b1;
	if(!_32) chunk_bits[15] = 1'b0;
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = 16'bxxxxxxxxxxxxxxxx;
	_RotateRight_data = chunk_bits;
end
always_comb begin // combinatorial _RotateRight_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_offset = 4'dx;
	_RotateRight_offset = chunk_offset;
end
endmodule

// RotateRight #(T: type bool #(), ARRAY_LEN: 16)
module RotateRight_T_type_bool_ARRAY_LEN_16(
	input clk,
	input wire[15:0] data,
	input wire[3:0] offset,
	output /*mux_wire*/ logic[15:0] rotated_data
);

/*mux_wire*/ logic[3:0] offset_bits;
/*mux_wire*/ logic[3:0] _UIntToBits_value;
wire[3:0] _UIntToBits_bits;
/*mux_wire*/ logic[15:0] rotate_stages[4:0];
/*mux_wire*/ logic[15:0] from;
wire[15:0] _3 = rotate_stages[0];
wire _4 = offset_bits[0];
wire _5 = from[15];
wire _6 = from[0];
wire _7 = offset_bits[0];
wire _8 = from[0];
wire _9 = from[1];
wire _10 = offset_bits[0];
wire _11 = from[1];
wire _12 = from[2];
wire _13 = offset_bits[0];
wire _14 = from[2];
wire _15 = from[3];
wire _16 = offset_bits[0];
wire _17 = from[3];
wire _18 = from[4];
wire _19 = offset_bits[0];
wire _20 = from[4];
wire _21 = from[5];
wire _22 = offset_bits[0];
wire _23 = from[5];
wire _24 = from[6];
wire _25 = offset_bits[0];
wire _26 = from[6];
wire _27 = from[7];
wire _28 = offset_bits[0];
wire _29 = from[7];
wire _30 = from[8];
wire _31 = offset_bits[0];
wire _32 = from[8];
wire _33 = from[9];
wire _34 = offset_bits[0];
wire _35 = from[9];
wire _36 = from[10];
wire _37 = offset_bits[0];
wire _38 = from[10];
wire _39 = from[11];
wire _40 = offset_bits[0];
wire _41 = from[11];
wire _42 = from[12];
wire _43 = offset_bits[0];
wire _44 = from[12];
wire _45 = from[13];
wire _46 = offset_bits[0];
wire _47 = from[13];
wire _48 = from[14];
wire _49 = offset_bits[0];
wire _50 = from[14];
wire _51 = from[15];
/*mux_wire*/ logic[15:0] from_2;
wire[15:0] _52 = rotate_stages[1];
wire _53 = offset_bits[1];
wire _54 = from_2[14];
wire _55 = from_2[0];
wire _56 = offset_bits[1];
wire _57 = from_2[15];
wire _58 = from_2[1];
wire _59 = offset_bits[1];
wire _60 = from_2[0];
wire _61 = from_2[2];
wire _62 = offset_bits[1];
wire _63 = from_2[1];
wire _64 = from_2[3];
wire _65 = offset_bits[1];
wire _66 = from_2[2];
wire _67 = from_2[4];
wire _68 = offset_bits[1];
wire _69 = from_2[3];
wire _70 = from_2[5];
wire _71 = offset_bits[1];
wire _72 = from_2[4];
wire _73 = from_2[6];
wire _74 = offset_bits[1];
wire _75 = from_2[5];
wire _76 = from_2[7];
wire _77 = offset_bits[1];
wire _78 = from_2[6];
wire _79 = from_2[8];
wire _80 = offset_bits[1];
wire _81 = from_2[7];
wire _82 = from_2[9];
wire _83 = offset_bits[1];
wire _84 = from_2[8];
wire _85 = from_2[10];
wire _86 = offset_bits[1];
wire _87 = from_2[9];
wire _88 = from_2[11];
wire _89 = offset_bits[1];
wire _90 = from_2[10];
wire _91 = from_2[12];
wire _92 = offset_bits[1];
wire _93 = from_2[11];
wire _94 = from_2[13];
wire _95 = offset_bits[1];
wire _96 = from_2[12];
wire _97 = from_2[14];
wire _98 = offset_bits[1];
wire _99 = from_2[13];
wire _100 = from_2[15];
/*mux_wire*/ logic[15:0] from_3;
wire[15:0] _101 = rotate_stages[2];
wire _102 = offset_bits[2];
wire _103 = from_3[12];
wire _104 = from_3[0];
wire _105 = offset_bits[2];
wire _106 = from_3[13];
wire _107 = from_3[1];
wire _108 = offset_bits[2];
wire _109 = from_3[14];
wire _110 = from_3[2];
wire _111 = offset_bits[2];
wire _112 = from_3[15];
wire _113 = from_3[3];
wire _114 = offset_bits[2];
wire _115 = from_3[0];
wire _116 = from_3[4];
wire _117 = offset_bits[2];
wire _118 = from_3[1];
wire _119 = from_3[5];
wire _120 = offset_bits[2];
wire _121 = from_3[2];
wire _122 = from_3[6];
wire _123 = offset_bits[2];
wire _124 = from_3[3];
wire _125 = from_3[7];
wire _126 = offset_bits[2];
wire _127 = from_3[4];
wire _128 = from_3[8];
wire _129 = offset_bits[2];
wire _130 = from_3[5];
wire _131 = from_3[9];
wire _132 = offset_bits[2];
wire _133 = from_3[6];
wire _134 = from_3[10];
wire _135 = offset_bits[2];
wire _136 = from_3[7];
wire _137 = from_3[11];
wire _138 = offset_bits[2];
wire _139 = from_3[8];
wire _140 = from_3[12];
wire _141 = offset_bits[2];
wire _142 = from_3[9];
wire _143 = from_3[13];
wire _144 = offset_bits[2];
wire _145 = from_3[10];
wire _146 = from_3[14];
wire _147 = offset_bits[2];
wire _148 = from_3[11];
wire _149 = from_3[15];
/*mux_wire*/ logic[15:0] from_4;
wire[15:0] _150 = rotate_stages[3];
wire _151 = offset_bits[3];
wire _152 = from_4[8];
wire _153 = from_4[0];
wire _154 = offset_bits[3];
wire _155 = from_4[9];
wire _156 = from_4[1];
wire _157 = offset_bits[3];
wire _158 = from_4[10];
wire _159 = from_4[2];
wire _160 = offset_bits[3];
wire _161 = from_4[11];
wire _162 = from_4[3];
wire _163 = offset_bits[3];
wire _164 = from_4[12];
wire _165 = from_4[4];
wire _166 = offset_bits[3];
wire _167 = from_4[13];
wire _168 = from_4[5];
wire _169 = offset_bits[3];
wire _170 = from_4[14];
wire _171 = from_4[6];
wire _172 = offset_bits[3];
wire _173 = from_4[15];
wire _174 = from_4[7];
wire _175 = offset_bits[3];
wire _176 = from_4[0];
wire _177 = from_4[8];
wire _178 = offset_bits[3];
wire _179 = from_4[1];
wire _180 = from_4[9];
wire _181 = offset_bits[3];
wire _182 = from_4[2];
wire _183 = from_4[10];
wire _184 = offset_bits[3];
wire _185 = from_4[3];
wire _186 = from_4[11];
wire _187 = offset_bits[3];
wire _188 = from_4[4];
wire _189 = from_4[12];
wire _190 = offset_bits[3];
wire _191 = from_4[5];
wire _192 = from_4[13];
wire _193 = offset_bits[3];
wire _194 = from_4[6];
wire _195 = from_4[14];
wire _196 = offset_bits[3];
wire _197 = from_4[7];
wire _198 = from_4[15];
wire[15:0] _199 = rotate_stages[4];
UIntToBits_NUM_BITS_4 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = 16'bxxxxxxxxxxxxxxxx;
	rotated_data = _199;
end
always_comb begin // combinatorial offset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	offset_bits = 4'bxxxx;
	offset_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 4'dx;
	_UIntToBits_value = offset;
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{16'bxxxxxxxxxxxxxxxx, 16'bxxxxxxxxxxxxxxxx, 16'bxxxxxxxxxxxxxxxx, 16'bxxxxxxxxxxxxxxxx, 16'bxxxxxxxxxxxxxxxx};
	rotate_stages[0] = data;
	if(_4) rotate_stages[1][0] = _5;
	if(!_4) rotate_stages[1][0] = _6;
	if(_7) rotate_stages[1][1] = _8;
	if(!_7) rotate_stages[1][1] = _9;
	if(_10) rotate_stages[1][2] = _11;
	if(!_10) rotate_stages[1][2] = _12;
	if(_13) rotate_stages[1][3] = _14;
	if(!_13) rotate_stages[1][3] = _15;
	if(_16) rotate_stages[1][4] = _17;
	if(!_16) rotate_stages[1][4] = _18;
	if(_19) rotate_stages[1][5] = _20;
	if(!_19) rotate_stages[1][5] = _21;
	if(_22) rotate_stages[1][6] = _23;
	if(!_22) rotate_stages[1][6] = _24;
	if(_25) rotate_stages[1][7] = _26;
	if(!_25) rotate_stages[1][7] = _27;
	if(_28) rotate_stages[1][8] = _29;
	if(!_28) rotate_stages[1][8] = _30;
	if(_31) rotate_stages[1][9] = _32;
	if(!_31) rotate_stages[1][9] = _33;
	if(_34) rotate_stages[1][10] = _35;
	if(!_34) rotate_stages[1][10] = _36;
	if(_37) rotate_stages[1][11] = _38;
	if(!_37) rotate_stages[1][11] = _39;
	if(_40) rotate_stages[1][12] = _41;
	if(!_40) rotate_stages[1][12] = _42;
	if(_43) rotate_stages[1][13] = _44;
	if(!_43) rotate_stages[1][13] = _45;
	if(_46) rotate_stages[1][14] = _47;
	if(!_46) rotate_stages[1][14] = _48;
	if(_49) rotate_stages[1][15] = _50;
	if(!_49) rotate_stages[1][15] = _51;
	if(_53) rotate_stages[2][0] = _54;
	if(!_53) rotate_stages[2][0] = _55;
	if(_56) rotate_stages[2][1] = _57;
	if(!_56) rotate_stages[2][1] = _58;
	if(_59) rotate_stages[2][2] = _60;
	if(!_59) rotate_stages[2][2] = _61;
	if(_62) rotate_stages[2][3] = _63;
	if(!_62) rotate_stages[2][3] = _64;
	if(_65) rotate_stages[2][4] = _66;
	if(!_65) rotate_stages[2][4] = _67;
	if(_68) rotate_stages[2][5] = _69;
	if(!_68) rotate_stages[2][5] = _70;
	if(_71) rotate_stages[2][6] = _72;
	if(!_71) rotate_stages[2][6] = _73;
	if(_74) rotate_stages[2][7] = _75;
	if(!_74) rotate_stages[2][7] = _76;
	if(_77) rotate_stages[2][8] = _78;
	if(!_77) rotate_stages[2][8] = _79;
	if(_80) rotate_stages[2][9] = _81;
	if(!_80) rotate_stages[2][9] = _82;
	if(_83) rotate_stages[2][10] = _84;
	if(!_83) rotate_stages[2][10] = _85;
	if(_86) rotate_stages[2][11] = _87;
	if(!_86) rotate_stages[2][11] = _88;
	if(_89) rotate_stages[2][12] = _90;
	if(!_89) rotate_stages[2][12] = _91;
	if(_92) rotate_stages[2][13] = _93;
	if(!_92) rotate_stages[2][13] = _94;
	if(_95) rotate_stages[2][14] = _96;
	if(!_95) rotate_stages[2][14] = _97;
	if(_98) rotate_stages[2][15] = _99;
	if(!_98) rotate_stages[2][15] = _100;
	if(_102) rotate_stages[3][0] = _103;
	if(!_102) rotate_stages[3][0] = _104;
	if(_105) rotate_stages[3][1] = _106;
	if(!_105) rotate_stages[3][1] = _107;
	if(_108) rotate_stages[3][2] = _109;
	if(!_108) rotate_stages[3][2] = _110;
	if(_111) rotate_stages[3][3] = _112;
	if(!_111) rotate_stages[3][3] = _113;
	if(_114) rotate_stages[3][4] = _115;
	if(!_114) rotate_stages[3][4] = _116;
	if(_117) rotate_stages[3][5] = _118;
	if(!_117) rotate_stages[3][5] = _119;
	if(_120) rotate_stages[3][6] = _121;
	if(!_120) rotate_stages[3][6] = _122;
	if(_123) rotate_stages[3][7] = _124;
	if(!_123) rotate_stages[3][7] = _125;
	if(_126) rotate_stages[3][8] = _127;
	if(!_126) rotate_stages[3][8] = _128;
	if(_129) rotate_stages[3][9] = _130;
	if(!_129) rotate_stages[3][9] = _131;
	if(_132) rotate_stages[3][10] = _133;
	if(!_132) rotate_stages[3][10] = _134;
	if(_135) rotate_stages[3][11] = _136;
	if(!_135) rotate_stages[3][11] = _137;
	if(_138) rotate_stages[3][12] = _139;
	if(!_138) rotate_stages[3][12] = _140;
	if(_141) rotate_stages[3][13] = _142;
	if(!_141) rotate_stages[3][13] = _143;
	if(_144) rotate_stages[3][14] = _145;
	if(!_144) rotate_stages[3][14] = _146;
	if(_147) rotate_stages[3][15] = _148;
	if(!_147) rotate_stages[3][15] = _149;
	if(_151) rotate_stages[4][0] = _152;
	if(!_151) rotate_stages[4][0] = _153;
	if(_154) rotate_stages[4][1] = _155;
	if(!_154) rotate_stages[4][1] = _156;
	if(_157) rotate_stages[4][2] = _158;
	if(!_157) rotate_stages[4][2] = _159;
	if(_160) rotate_stages[4][3] = _161;
	if(!_160) rotate_stages[4][3] = _162;
	if(_163) rotate_stages[4][4] = _164;
	if(!_163) rotate_stages[4][4] = _165;
	if(_166) rotate_stages[4][5] = _167;
	if(!_166) rotate_stages[4][5] = _168;
	if(_169) rotate_stages[4][6] = _170;
	if(!_169) rotate_stages[4][6] = _171;
	if(_172) rotate_stages[4][7] = _173;
	if(!_172) rotate_stages[4][7] = _174;
	if(_175) rotate_stages[4][8] = _176;
	if(!_175) rotate_stages[4][8] = _177;
	if(_178) rotate_stages[4][9] = _179;
	if(!_178) rotate_stages[4][9] = _180;
	if(_181) rotate_stages[4][10] = _182;
	if(!_181) rotate_stages[4][10] = _183;
	if(_184) rotate_stages[4][11] = _185;
	if(!_184) rotate_stages[4][11] = _186;
	if(_187) rotate_stages[4][12] = _188;
	if(!_187) rotate_stages[4][12] = _189;
	if(_190) rotate_stages[4][13] = _191;
	if(!_190) rotate_stages[4][13] = _192;
	if(_193) rotate_stages[4][14] = _194;
	if(!_193) rotate_stages[4][14] = _195;
	if(_196) rotate_stages[4][15] = _197;
	if(!_196) rotate_stages[4][15] = _198;
end
always_comb begin // combinatorial from
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from = 16'bxxxxxxxxxxxxxxxx;
	from = _3;
end
always_comb begin // combinatorial from_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_2 = 16'bxxxxxxxxxxxxxxxx;
	from_2 = _52;
end
always_comb begin // combinatorial from_3
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_3 = 16'bxxxxxxxxxxxxxxxx;
	from_3 = _101;
end
always_comb begin // combinatorial from_4
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_4 = 16'bxxxxxxxxxxxxxxxx;
	from_4 = _150;
end
endmodule

// RotateRight #(T: type bool #()[32], ARRAY_LEN: 16)
module RotateRight_T_type_bool_32_ARRAY_LEN_16(
	input clk,
	input wire[31:0] data[15:0],
	input wire[3:0] offset,
	output /*mux_wire*/ logic[31:0] rotated_data[15:0]
);

genvar _g0;
/*mux_wire*/ logic[3:0] offset_bits;
/*mux_wire*/ logic[3:0] _UIntToBits_value;
wire[3:0] _UIntToBits_bits;
/*mux_wire*/ logic[31:0] rotate_stages[4:0][15:0];
/*mux_wire*/ logic[31:0] from[15:0];
wire[31:0] _3[15:0];
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _3[_g0] = rotate_stages[0][_g0];
end
endgenerate
wire _4 = offset_bits[0];
wire[31:0] _5 = from[15];
wire[31:0] _6 = from[0];
wire _7 = offset_bits[0];
wire[31:0] _8 = from[0];
wire[31:0] _9 = from[1];
wire _10 = offset_bits[0];
wire[31:0] _11 = from[1];
wire[31:0] _12 = from[2];
wire _13 = offset_bits[0];
wire[31:0] _14 = from[2];
wire[31:0] _15 = from[3];
wire _16 = offset_bits[0];
wire[31:0] _17 = from[3];
wire[31:0] _18 = from[4];
wire _19 = offset_bits[0];
wire[31:0] _20 = from[4];
wire[31:0] _21 = from[5];
wire _22 = offset_bits[0];
wire[31:0] _23 = from[5];
wire[31:0] _24 = from[6];
wire _25 = offset_bits[0];
wire[31:0] _26 = from[6];
wire[31:0] _27 = from[7];
wire _28 = offset_bits[0];
wire[31:0] _29 = from[7];
wire[31:0] _30 = from[8];
wire _31 = offset_bits[0];
wire[31:0] _32 = from[8];
wire[31:0] _33 = from[9];
wire _34 = offset_bits[0];
wire[31:0] _35 = from[9];
wire[31:0] _36 = from[10];
wire _37 = offset_bits[0];
wire[31:0] _38 = from[10];
wire[31:0] _39 = from[11];
wire _40 = offset_bits[0];
wire[31:0] _41 = from[11];
wire[31:0] _42 = from[12];
wire _43 = offset_bits[0];
wire[31:0] _44 = from[12];
wire[31:0] _45 = from[13];
wire _46 = offset_bits[0];
wire[31:0] _47 = from[13];
wire[31:0] _48 = from[14];
wire _49 = offset_bits[0];
wire[31:0] _50 = from[14];
wire[31:0] _51 = from[15];
/*mux_wire*/ logic[31:0] from_2[15:0];
wire[31:0] _52[15:0];
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _52[_g0] = rotate_stages[1][_g0];
end
endgenerate
wire _53 = offset_bits[1];
wire[31:0] _54 = from_2[14];
wire[31:0] _55 = from_2[0];
wire _56 = offset_bits[1];
wire[31:0] _57 = from_2[15];
wire[31:0] _58 = from_2[1];
wire _59 = offset_bits[1];
wire[31:0] _60 = from_2[0];
wire[31:0] _61 = from_2[2];
wire _62 = offset_bits[1];
wire[31:0] _63 = from_2[1];
wire[31:0] _64 = from_2[3];
wire _65 = offset_bits[1];
wire[31:0] _66 = from_2[2];
wire[31:0] _67 = from_2[4];
wire _68 = offset_bits[1];
wire[31:0] _69 = from_2[3];
wire[31:0] _70 = from_2[5];
wire _71 = offset_bits[1];
wire[31:0] _72 = from_2[4];
wire[31:0] _73 = from_2[6];
wire _74 = offset_bits[1];
wire[31:0] _75 = from_2[5];
wire[31:0] _76 = from_2[7];
wire _77 = offset_bits[1];
wire[31:0] _78 = from_2[6];
wire[31:0] _79 = from_2[8];
wire _80 = offset_bits[1];
wire[31:0] _81 = from_2[7];
wire[31:0] _82 = from_2[9];
wire _83 = offset_bits[1];
wire[31:0] _84 = from_2[8];
wire[31:0] _85 = from_2[10];
wire _86 = offset_bits[1];
wire[31:0] _87 = from_2[9];
wire[31:0] _88 = from_2[11];
wire _89 = offset_bits[1];
wire[31:0] _90 = from_2[10];
wire[31:0] _91 = from_2[12];
wire _92 = offset_bits[1];
wire[31:0] _93 = from_2[11];
wire[31:0] _94 = from_2[13];
wire _95 = offset_bits[1];
wire[31:0] _96 = from_2[12];
wire[31:0] _97 = from_2[14];
wire _98 = offset_bits[1];
wire[31:0] _99 = from_2[13];
wire[31:0] _100 = from_2[15];
/*mux_wire*/ logic[31:0] from_3[15:0];
wire[31:0] _101[15:0];
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _101[_g0] = rotate_stages[2][_g0];
end
endgenerate
wire _102 = offset_bits[2];
wire[31:0] _103 = from_3[12];
wire[31:0] _104 = from_3[0];
wire _105 = offset_bits[2];
wire[31:0] _106 = from_3[13];
wire[31:0] _107 = from_3[1];
wire _108 = offset_bits[2];
wire[31:0] _109 = from_3[14];
wire[31:0] _110 = from_3[2];
wire _111 = offset_bits[2];
wire[31:0] _112 = from_3[15];
wire[31:0] _113 = from_3[3];
wire _114 = offset_bits[2];
wire[31:0] _115 = from_3[0];
wire[31:0] _116 = from_3[4];
wire _117 = offset_bits[2];
wire[31:0] _118 = from_3[1];
wire[31:0] _119 = from_3[5];
wire _120 = offset_bits[2];
wire[31:0] _121 = from_3[2];
wire[31:0] _122 = from_3[6];
wire _123 = offset_bits[2];
wire[31:0] _124 = from_3[3];
wire[31:0] _125 = from_3[7];
wire _126 = offset_bits[2];
wire[31:0] _127 = from_3[4];
wire[31:0] _128 = from_3[8];
wire _129 = offset_bits[2];
wire[31:0] _130 = from_3[5];
wire[31:0] _131 = from_3[9];
wire _132 = offset_bits[2];
wire[31:0] _133 = from_3[6];
wire[31:0] _134 = from_3[10];
wire _135 = offset_bits[2];
wire[31:0] _136 = from_3[7];
wire[31:0] _137 = from_3[11];
wire _138 = offset_bits[2];
wire[31:0] _139 = from_3[8];
wire[31:0] _140 = from_3[12];
wire _141 = offset_bits[2];
wire[31:0] _142 = from_3[9];
wire[31:0] _143 = from_3[13];
wire _144 = offset_bits[2];
wire[31:0] _145 = from_3[10];
wire[31:0] _146 = from_3[14];
wire _147 = offset_bits[2];
wire[31:0] _148 = from_3[11];
wire[31:0] _149 = from_3[15];
/*mux_wire*/ logic[31:0] from_4[15:0];
wire[31:0] _150[15:0];
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _150[_g0] = rotate_stages[3][_g0];
end
endgenerate
wire _151 = offset_bits[3];
wire[31:0] _152 = from_4[8];
wire[31:0] _153 = from_4[0];
wire _154 = offset_bits[3];
wire[31:0] _155 = from_4[9];
wire[31:0] _156 = from_4[1];
wire _157 = offset_bits[3];
wire[31:0] _158 = from_4[10];
wire[31:0] _159 = from_4[2];
wire _160 = offset_bits[3];
wire[31:0] _161 = from_4[11];
wire[31:0] _162 = from_4[3];
wire _163 = offset_bits[3];
wire[31:0] _164 = from_4[12];
wire[31:0] _165 = from_4[4];
wire _166 = offset_bits[3];
wire[31:0] _167 = from_4[13];
wire[31:0] _168 = from_4[5];
wire _169 = offset_bits[3];
wire[31:0] _170 = from_4[14];
wire[31:0] _171 = from_4[6];
wire _172 = offset_bits[3];
wire[31:0] _173 = from_4[15];
wire[31:0] _174 = from_4[7];
wire _175 = offset_bits[3];
wire[31:0] _176 = from_4[0];
wire[31:0] _177 = from_4[8];
wire _178 = offset_bits[3];
wire[31:0] _179 = from_4[1];
wire[31:0] _180 = from_4[9];
wire _181 = offset_bits[3];
wire[31:0] _182 = from_4[2];
wire[31:0] _183 = from_4[10];
wire _184 = offset_bits[3];
wire[31:0] _185 = from_4[3];
wire[31:0] _186 = from_4[11];
wire _187 = offset_bits[3];
wire[31:0] _188 = from_4[4];
wire[31:0] _189 = from_4[12];
wire _190 = offset_bits[3];
wire[31:0] _191 = from_4[5];
wire[31:0] _192 = from_4[13];
wire _193 = offset_bits[3];
wire[31:0] _194 = from_4[6];
wire[31:0] _195 = from_4[14];
wire _196 = offset_bits[3];
wire[31:0] _197 = from_4[7];
wire[31:0] _198 = from_4[15];
wire[31:0] _199[15:0];
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _199[_g0] = rotate_stages[4][_g0];
end
endgenerate
UIntToBits_NUM_BITS_4 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
rotated_data[_v0] = _199[_v0];
end
end
always_comb begin // combinatorial offset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	offset_bits = 4'bxxxx;
	offset_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 4'dx;
	_UIntToBits_value = offset;
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{'{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
rotate_stages[0][_v0] = data[_v0];
end
	if(_4) rotate_stages[1][0] = _5;
	if(!_4) rotate_stages[1][0] = _6;
	if(_7) rotate_stages[1][1] = _8;
	if(!_7) rotate_stages[1][1] = _9;
	if(_10) rotate_stages[1][2] = _11;
	if(!_10) rotate_stages[1][2] = _12;
	if(_13) rotate_stages[1][3] = _14;
	if(!_13) rotate_stages[1][3] = _15;
	if(_16) rotate_stages[1][4] = _17;
	if(!_16) rotate_stages[1][4] = _18;
	if(_19) rotate_stages[1][5] = _20;
	if(!_19) rotate_stages[1][5] = _21;
	if(_22) rotate_stages[1][6] = _23;
	if(!_22) rotate_stages[1][6] = _24;
	if(_25) rotate_stages[1][7] = _26;
	if(!_25) rotate_stages[1][7] = _27;
	if(_28) rotate_stages[1][8] = _29;
	if(!_28) rotate_stages[1][8] = _30;
	if(_31) rotate_stages[1][9] = _32;
	if(!_31) rotate_stages[1][9] = _33;
	if(_34) rotate_stages[1][10] = _35;
	if(!_34) rotate_stages[1][10] = _36;
	if(_37) rotate_stages[1][11] = _38;
	if(!_37) rotate_stages[1][11] = _39;
	if(_40) rotate_stages[1][12] = _41;
	if(!_40) rotate_stages[1][12] = _42;
	if(_43) rotate_stages[1][13] = _44;
	if(!_43) rotate_stages[1][13] = _45;
	if(_46) rotate_stages[1][14] = _47;
	if(!_46) rotate_stages[1][14] = _48;
	if(_49) rotate_stages[1][15] = _50;
	if(!_49) rotate_stages[1][15] = _51;
	if(_53) rotate_stages[2][0] = _54;
	if(!_53) rotate_stages[2][0] = _55;
	if(_56) rotate_stages[2][1] = _57;
	if(!_56) rotate_stages[2][1] = _58;
	if(_59) rotate_stages[2][2] = _60;
	if(!_59) rotate_stages[2][2] = _61;
	if(_62) rotate_stages[2][3] = _63;
	if(!_62) rotate_stages[2][3] = _64;
	if(_65) rotate_stages[2][4] = _66;
	if(!_65) rotate_stages[2][4] = _67;
	if(_68) rotate_stages[2][5] = _69;
	if(!_68) rotate_stages[2][5] = _70;
	if(_71) rotate_stages[2][6] = _72;
	if(!_71) rotate_stages[2][6] = _73;
	if(_74) rotate_stages[2][7] = _75;
	if(!_74) rotate_stages[2][7] = _76;
	if(_77) rotate_stages[2][8] = _78;
	if(!_77) rotate_stages[2][8] = _79;
	if(_80) rotate_stages[2][9] = _81;
	if(!_80) rotate_stages[2][9] = _82;
	if(_83) rotate_stages[2][10] = _84;
	if(!_83) rotate_stages[2][10] = _85;
	if(_86) rotate_stages[2][11] = _87;
	if(!_86) rotate_stages[2][11] = _88;
	if(_89) rotate_stages[2][12] = _90;
	if(!_89) rotate_stages[2][12] = _91;
	if(_92) rotate_stages[2][13] = _93;
	if(!_92) rotate_stages[2][13] = _94;
	if(_95) rotate_stages[2][14] = _96;
	if(!_95) rotate_stages[2][14] = _97;
	if(_98) rotate_stages[2][15] = _99;
	if(!_98) rotate_stages[2][15] = _100;
	if(_102) rotate_stages[3][0] = _103;
	if(!_102) rotate_stages[3][0] = _104;
	if(_105) rotate_stages[3][1] = _106;
	if(!_105) rotate_stages[3][1] = _107;
	if(_108) rotate_stages[3][2] = _109;
	if(!_108) rotate_stages[3][2] = _110;
	if(_111) rotate_stages[3][3] = _112;
	if(!_111) rotate_stages[3][3] = _113;
	if(_114) rotate_stages[3][4] = _115;
	if(!_114) rotate_stages[3][4] = _116;
	if(_117) rotate_stages[3][5] = _118;
	if(!_117) rotate_stages[3][5] = _119;
	if(_120) rotate_stages[3][6] = _121;
	if(!_120) rotate_stages[3][6] = _122;
	if(_123) rotate_stages[3][7] = _124;
	if(!_123) rotate_stages[3][7] = _125;
	if(_126) rotate_stages[3][8] = _127;
	if(!_126) rotate_stages[3][8] = _128;
	if(_129) rotate_stages[3][9] = _130;
	if(!_129) rotate_stages[3][9] = _131;
	if(_132) rotate_stages[3][10] = _133;
	if(!_132) rotate_stages[3][10] = _134;
	if(_135) rotate_stages[3][11] = _136;
	if(!_135) rotate_stages[3][11] = _137;
	if(_138) rotate_stages[3][12] = _139;
	if(!_138) rotate_stages[3][12] = _140;
	if(_141) rotate_stages[3][13] = _142;
	if(!_141) rotate_stages[3][13] = _143;
	if(_144) rotate_stages[3][14] = _145;
	if(!_144) rotate_stages[3][14] = _146;
	if(_147) rotate_stages[3][15] = _148;
	if(!_147) rotate_stages[3][15] = _149;
	if(_151) rotate_stages[4][0] = _152;
	if(!_151) rotate_stages[4][0] = _153;
	if(_154) rotate_stages[4][1] = _155;
	if(!_154) rotate_stages[4][1] = _156;
	if(_157) rotate_stages[4][2] = _158;
	if(!_157) rotate_stages[4][2] = _159;
	if(_160) rotate_stages[4][3] = _161;
	if(!_160) rotate_stages[4][3] = _162;
	if(_163) rotate_stages[4][4] = _164;
	if(!_163) rotate_stages[4][4] = _165;
	if(_166) rotate_stages[4][5] = _167;
	if(!_166) rotate_stages[4][5] = _168;
	if(_169) rotate_stages[4][6] = _170;
	if(!_169) rotate_stages[4][6] = _171;
	if(_172) rotate_stages[4][7] = _173;
	if(!_172) rotate_stages[4][7] = _174;
	if(_175) rotate_stages[4][8] = _176;
	if(!_175) rotate_stages[4][8] = _177;
	if(_178) rotate_stages[4][9] = _179;
	if(!_178) rotate_stages[4][9] = _180;
	if(_181) rotate_stages[4][10] = _182;
	if(!_181) rotate_stages[4][10] = _183;
	if(_184) rotate_stages[4][11] = _185;
	if(!_184) rotate_stages[4][11] = _186;
	if(_187) rotate_stages[4][12] = _188;
	if(!_187) rotate_stages[4][12] = _189;
	if(_190) rotate_stages[4][13] = _191;
	if(!_190) rotate_stages[4][13] = _192;
	if(_193) rotate_stages[4][14] = _194;
	if(!_193) rotate_stages[4][14] = _195;
	if(_196) rotate_stages[4][15] = _197;
	if(!_196) rotate_stages[4][15] = _198;
end
always_comb begin // combinatorial from
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
from[_v0] = _3[_v0];
end
end
always_comb begin // combinatorial from_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_2 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
from_2[_v0] = _52[_v0];
end
end
always_comb begin // combinatorial from_3
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_3 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
from_3[_v0] = _101[_v0];
end
end
always_comb begin // combinatorial from_4
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_4 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
from_4[_v0] = _150[_v0];
end
end
endmodule

// axi_array_burst_reader #(AXI_WIDTH: 512, ADDR_ALIGN: 4, COUNT_TO: 68719476736, ATO: 18446744073709551616)
module axi_array_burst_reader_AXI_WIDTH_512_ADDR_ALIGN_4_COUNT_TO_68719476736_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*state*/ logic arvalid,
	input wire arready,
	output /*state*/ logic[63:0] araddr,
	output /*state*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[511:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic element_packet_valid,
	output /*mux_wire*/ logic[31:0] elements[15:0],
	output /*mux_wire*/ logic[3:0] chunk_offset,
	output /*mux_wire*/ logic[4:0] chunk_length,
	output /*mux_wire*/ logic last,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[35:0] count
);

/*latency*/ logic _arvalid_D1; always_ff @(posedge aclk) begin _arvalid_D1 <= arvalid; end
/*latency*/ logic _request_new_burst_D1; always_ff @(posedge aclk) begin _request_new_burst_D1 <= request_new_burst; end
genvar _g0;
localparam[1:0] _1 = 2'b01;
localparam[2:0] _2 = 3'b000;
localparam[3:0] _3 = 4'b0010;
/*mux_wire*/ logic[1:0] _rresp;
/*mux_wire*/ logic _rlast;
/*state*/ logic[11:0] num_in_flight;
/*state*/ logic last_burst_in_flight;
/*mux_wire*/ logic[63:0] next_araddr;
/*latency*/ logic[63:0] _next_araddr_D0; always_ff @(posedge aclk) begin _next_araddr_D0 <= next_araddr; end
wire[57:0] _cur_start_chunk_addr_old;
/*mux_wire*/ logic[57:0] _BitwiseIntConcat_upper;
/*mux_wire*/ logic[5:0] _BitwiseIntConcat_lower;
wire[63:0] _BitwiseIntConcat_v;
/*mux_wire*/ logic[5:0] next_arlen;
/*mux_wire*/ logic next_last_burst_in_flight;
/*latency*/ logic _next_last_burst_in_flight_D0; always_ff @(posedge aclk) begin _next_last_burst_in_flight_D0 <= next_last_burst_in_flight; end
/*mux_wire*/ logic[51:0] cur_burst_addr;
/*mux_wire*/ logic[5:0] cur_align;
/*mux_wire*/ logic[57:0] _BitwiseIntSplit_v;
wire[51:0] _BitwiseIntSplit_upper;
wire[5:0] _BitwiseIntSplit_lower;
/*mux_wire*/ logic chunks_are_left;
/*latency*/ logic _chunks_are_left_D0; always_ff @(posedge aclk) begin _chunks_are_left_D0 <= chunks_are_left; end
wire[32:0] _num_chunks_left_old;
/*latency*/ logic[32:0] __num_chunks_left_old_N1; always_ff @(posedge aclk) begin __num_chunks_left_old_N1 <= _num_chunks_left_old; end
/*latency*/ logic[32:0] __num_chunks_left_old_D0; always_ff @(posedge aclk) begin __num_chunks_left_old_D0 <= __num_chunks_left_old_N1; end
wire _14;
assign _14 = _num_chunks_left_old > 1'd0;
/*latency*/ logic __14_N1; always_ff @(posedge aclk) begin __14_N1 <= _14; end
/*mux_wire*/ logic[5:0] max_chunks_in_this_burst;
/*latency*/ logic[5:0] _max_chunks_in_this_burst_D0; always_ff @(posedge aclk) begin _max_chunks_in_this_burst_D0 <= max_chunks_in_this_burst; end
wire[5:0] _18;
assign _18 = 6'd63 - cur_align;
wire[6:0] _22;
assign _22 = max_chunks_in_this_burst + 1'd1;
wire _23;
assign _23 = __num_chunks_left_old_N1 <= _22;
/*latency*/ logic __23_D0; always_ff @(posedge aclk) begin __23_D0 <= _23; end
/*mux_wire*/ logic[32:0] _IntNarrow_in;
wire[6:0] _IntNarrow_out;
wire[5:0] _26;
assign _26 = _IntNarrow_out - 1'd1;
/*latency*/ logic[5:0] __26_D0; always_ff @(posedge aclk) begin __26_D0 <= _26; end
/*mux_wire*/ logic may_next_arvalid;
/*latency*/ logic _may_next_arvalid_D1; always_ff @(posedge aclk) begin _may_next_arvalid_D1 <= may_next_arvalid; end
wire _num_chunks_left_may_update;
wire _30;
assign _30 = _chunks_are_left_D0 & _num_chunks_left_may_update;
wire _cur_start_chunk_addr_may_update;
wire _32;
assign _32 = _30 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
wire _34;
assign _34 = _32 & _LatencyOffset_out;
wire signed[11:0] _37;
assign _37 = max_in_flight - 7'd64;
wire _38;
assign _38 = $signed({1'b0, num_in_flight}) <= _37;
wire _39;
assign _39 = _34 & _38;
/*mux_wire*/ logic[52:0] next_burst_addr;
wire[52:0] _45;
assign _45 = cur_burst_addr + 1'd1;
/*latency*/ logic[52:0] __45_D0; always_ff @(posedge aclk) begin __45_D0 <= _45; end
/*latency*/ logic[52:0] __45_D1; always_ff @(posedge aclk) begin __45_D1 <= __45_D0; end
/*mux_wire*/ logic[52:0] _BitwiseIntConcat_2_upper;
/*mux_wire*/ logic[5:0] _BitwiseIntConcat_2_lower;
wire[58:0] _BitwiseIntConcat_2_v;
/*mux_wire*/ logic[58:0] _IntNarrow_2_in;
wire[57:0] _IntNarrow_2_out;
/*mux_wire*/ logic _cur_start_chunk_addr_update;
/*mux_wire*/ logic[57:0] _cur_start_chunk_addr_new;
/*mux_wire*/ logic[32:0] next_num_chunks_left;
wire[6:0] _53;
assign _53 = next_arlen + 1'd1;
wire signed[33:0] _54;
assign _54 = __num_chunks_left_old_D0 - _53;
/*mux_wire*/ logic signed[33:0] _IntNarrow_3_in;
wire[32:0] _IntNarrow_3_out;
/*mux_wire*/ logic _num_chunks_left_update;
/*mux_wire*/ logic[32:0] _num_chunks_left_new;
/*mux_wire*/ logic _BoolToInt_i;
wire[0:0] _BoolToInt_o;
wire signed[12:0] _64;
assign _64 = num_in_flight - _BoolToInt_o;
wire _66;
assign _66 = !arvalid;
wire _68;
assign _68 = _66 & may_next_arvalid;
wire[6:0] _71;
assign _71 = next_arlen + 1'd1;
/*mux_wire*/ logic _Ternary_cond;
/*mux_wire*/ logic[6:0] _Ternary_a;
/*mux_wire*/ logic[6:0] _Ternary_b;
wire[6:0] _Ternary_o;
wire signed[12:0] _73;
assign _73 = _64 + $signed({1'b0, _Ternary_o});
/*mux_wire*/ logic signed[12:0] _IntNarrow_4_in;
wire[11:0] _IntNarrow_4_out;
/*state*/ logic[4:0] final_chunk_align;
/*state*/ logic[3:0] cur_chunk_align;
/*mux_wire*/ logic[31:0] elements_2[15:0];
wire[31:0] _75;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _75[_g0] = rdata[_g0];
end
endgenerate
wire[31:0] _76;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _76[_g0] = rdata[32 + _g0];
end
endgenerate
wire[31:0] _77;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _77[_g0] = rdata[64 + _g0];
end
endgenerate
wire[31:0] _78;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _78[_g0] = rdata[96 + _g0];
end
endgenerate
wire[31:0] _79;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _79[_g0] = rdata[128 + _g0];
end
endgenerate
wire[31:0] _80;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _80[_g0] = rdata[160 + _g0];
end
endgenerate
wire[31:0] _81;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _81[_g0] = rdata[192 + _g0];
end
endgenerate
wire[31:0] _82;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _82[_g0] = rdata[224 + _g0];
end
endgenerate
wire[31:0] _83;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _83[_g0] = rdata[256 + _g0];
end
endgenerate
wire[31:0] _84;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _84[_g0] = rdata[288 + _g0];
end
endgenerate
wire[31:0] _85;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _85[_g0] = rdata[320 + _g0];
end
endgenerate
wire[31:0] _86;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _86[_g0] = rdata[352 + _g0];
end
endgenerate
wire[31:0] _87;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _87[_g0] = rdata[384 + _g0];
end
endgenerate
wire[31:0] _88;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _88[_g0] = rdata[416 + _g0];
end
endgenerate
wire[31:0] _89;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _89[_g0] = rdata[448 + _g0];
end
endgenerate
wire[31:0] _90;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _90[_g0] = rdata[480 + _g0];
end
endgenerate
/*mux_wire*/ logic[4:0] num_chunk_elements;
/*mux_wire*/ logic is_last;
wire _93;
assign _93 = num_in_flight == 1'd1;
wire _95;
assign _95 = _93 & last_burst_in_flight;
wire signed[5:0] _99;
assign _99 = final_chunk_align - cur_chunk_align;
/*mux_wire*/ logic signed[5:0] _IntNarrow_5_in;
wire[4:0] _IntNarrow_5_out;
wire[4:0] _101;
assign _101 = 5'd16 - cur_chunk_align;
wire _109;
assign _109 = !chunks_are_left;
/*latency*/ logic __109_D0; always_ff @(posedge aclk) begin __109_D0 <= _109; end
wire _111;
assign _111 = __109_D0 & _num_chunks_left_may_update;
wire _113;
assign _113 = _111 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic[57:0] chunk_addr;
/*latency*/ logic[57:0] _chunk_addr_D1; always_ff @(posedge aclk) begin _chunk_addr_D1 <= chunk_addr; end
/*mux_wire*/ logic[3:0] element_in_chunk_align;
wire[61:0] _115;
assign _115 = start_addr / 3'd4;
/*mux_wire*/ logic[61:0] _BitwiseIntSplit_2_v;
wire[57:0] _BitwiseIntSplit_2_upper;
wire[3:0] _BitwiseIntSplit_2_lower;
/*mux_wire*/ logic[32:0] chunk_count_bits;
/*mux_wire*/ logic[3:0] final_alignment;
wire[36:0] _118;
assign _118 = count + element_in_chunk_align;
/*mux_wire*/ logic[36:0] _BitwiseIntSplit_3_v;
wire[32:0] _BitwiseIntSplit_3_upper;
wire[3:0] _BitwiseIntSplit_3_lower;
/*mux_wire*/ logic[32:0] num_chunks;
/*mux_wire*/ logic is_no_chunks;
wire _121;
assign _121 = chunk_count_bits == 1'd0;
wire _127;
assign _127 = final_alignment != 1'd0;
/*mux_wire*/ logic _BoolToInt_2_i;
wire[0:0] _BoolToInt_2_o;
wire[32:0] _128;
assign _128 = chunk_count_bits + _BoolToInt_2_o;
wire _134;
assign _134 = !is_no_chunks;
wire _137;
assign _137 = final_alignment == 1'd0;
wire _138;
assign _138 = _134 & _137;
/*mux_wire*/ logic _BoolToInt_3_i;
wire[0:0] _BoolToInt_3_o;
/*mux_wire*/ logic[0:0] _BitwiseIntConcat_3_upper;
/*mux_wire*/ logic[3:0] _BitwiseIntConcat_3_lower;
wire[4:0] _BitwiseIntConcat_3_v;
wire _142;
assign _142 = !aresetn;
/*mux_wire*/ logic _cur_start_chunk_addr_rst;
wire _144;
assign _144 = !aresetn;
/*mux_wire*/ logic _num_chunks_left_rst;
wire _146;
assign _146 = !aresetn;
SlowState_T_type_int_FROM_0_TO_288230376151711744_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1 cur_start_chunk_addr(
	.clk(aclk),
	.rst(_cur_start_chunk_addr_rst),
	.old(_cur_start_chunk_addr_old),
	.may_update(_cur_start_chunk_addr_may_update),
	.update(_cur_start_chunk_addr_update),
	.new_1(_cur_start_chunk_addr_new)
);
SlowState_T_type_int_FROM_0_TO_4294967299_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0 num_chunks_left(
	.clk(aclk),
	.rst(_num_chunks_left_rst),
	.old(_num_chunks_left_old),
	.may_update(_num_chunks_left_may_update),
	.update(_num_chunks_left_update),
	.new_1(_num_chunks_left_new)
);
BitwiseIntConcat_UPPER_TO_288230376151711744_LOWER_BITS_6 BitwiseIntConcat(
	.clk(aclk),
	.upper(_BitwiseIntConcat_upper),
	.lower(_BitwiseIntConcat_lower),
	.v(_BitwiseIntConcat_v)
);
BitwiseIntSplit_TO_288230376151711744_LOWER_BITS_6 BitwiseIntSplit(
	.clk(aclk),
	.v(_BitwiseIntSplit_v),
	.upper(_BitwiseIntSplit_upper),
	.lower(_BitwiseIntSplit_lower)
);
IntNarrow_FROM_I_0_TO_I_4294967299_FROM_1_TO_65 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
LatencyOffset_T_type_bool_OFFSET_192 LatencyOffset(
	.clk(aclk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
BitwiseIntConcat_UPPER_TO_4503599627370497_LOWER_BITS_6 BitwiseIntConcat_2(
	.clk(aclk),
	.upper(_BitwiseIntConcat_2_upper),
	.lower(_BitwiseIntConcat_2_lower),
	.v(_BitwiseIntConcat_2_v)
);
IntNarrow_FROM_I_0_TO_I_288230376151711808_FROM_0_TO_288230376151711744 IntNarrow_2(
	.clk(aclk),
	.in(_IntNarrow_2_in),
	.out(_IntNarrow_2_out)
);
IntNarrow_FROM_I_64_TO_I_4294967298_FROM_0_TO_4294967299 IntNarrow_3(
	.clk(aclk),
	.in(_IntNarrow_3_in),
	.out(_IntNarrow_3_out)
);
BoolToInt BoolToInt(
	.clk(aclk),
	.i(_BoolToInt_i),
	.o(_BoolToInt_o)
);
Ternary_T_type_int_FROM_0_TO_65 Ternary(
	.clk(aclk),
	.cond(_Ternary_cond),
	.a(_Ternary_a),
	.b(_Ternary_b),
	.o(_Ternary_o)
);
IntNarrow_FROM_I_1_TO_I_3256_FROM_0_TO_3192 IntNarrow_4(
	.clk(aclk),
	.in(_IntNarrow_4_in),
	.out(_IntNarrow_4_out)
);
IntNarrow_FROM_I_15_TO_I_32_FROM_0_TO_17 IntNarrow_5(
	.clk(aclk),
	.in(_IntNarrow_5_in),
	.out(_IntNarrow_5_out)
);
BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_4 BitwiseIntSplit_2(
	.clk(aclk),
	.v(_BitwiseIntSplit_2_v),
	.upper(_BitwiseIntSplit_2_upper),
	.lower(_BitwiseIntSplit_2_lower)
);
BitwiseIntSplit_TO_68719476751_LOWER_BITS_4 BitwiseIntSplit_3(
	.clk(aclk),
	.v(_BitwiseIntSplit_3_v),
	.upper(_BitwiseIntSplit_3_upper),
	.lower(_BitwiseIntSplit_3_lower)
);
BoolToInt BoolToInt_2(
	.clk(aclk),
	.i(_BoolToInt_2_i),
	.o(_BoolToInt_2_o)
);
BoolToInt BoolToInt_3(
	.clk(aclk),
	.i(_BoolToInt_3_i),
	.o(_BoolToInt_3_o)
);
BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_4 BitwiseIntConcat_3(
	.clk(aclk),
	.upper(_BitwiseIntConcat_3_upper),
	.lower(_BitwiseIntConcat_3_lower),
	.v(_BitwiseIntConcat_3_v)
);
always_ff @(posedge aclk) begin // state arvalid
	if(arvalid) if(arready) arvalid <= 1'b0;
	if(!arvalid) if(may_next_arvalid) arvalid <= 1'b1;
	if(_146) arvalid <= 1'b0;
end
always_ff @(posedge aclk) begin // state araddr
	if(!arvalid) if(may_next_arvalid) araddr <= _next_araddr_D0;
end
always_ff @(posedge aclk) begin // state arlen
	if(!arvalid) if(may_next_arvalid) arlen <= next_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = 3'd6;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _1;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _2;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _3;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = 1'd0;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = 1'd0;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rresp = 2'bxx;
	_rresp = rresp;
end
always_comb begin // combinatorial _rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rlast = 1'bx;
	_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_rlast = _rlast;
end
always_comb begin // combinatorial element_packet_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_packet_valid = 1'bx;
	element_packet_valid = 1'b0;
	if(rvalid) element_packet_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	element_packet_valid = element_packet_valid;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
if(rvalid) elements[_v0] = elements_2[_v0];
end
end
always_comb begin // combinatorial chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_offset = 4'dx;
	if(rvalid) chunk_offset = cur_chunk_align;
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 5'dx;
	if(rvalid) chunk_length = num_chunk_elements;
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(rvalid) last = is_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state num_in_flight
	num_in_flight <= _IntNarrow_4_out;
	if(_146) num_in_flight <= 1'd0;
end
always_ff @(posedge aclk) begin // state last_burst_in_flight
	if(!arvalid) if(may_next_arvalid) last_burst_in_flight <= _next_last_burst_in_flight_D0;
end
always_comb begin // combinatorial next_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_araddr = 64'dx;
	next_araddr = _BitwiseIntConcat_v;
end
always_comb begin // combinatorial _BitwiseIntConcat_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_upper = 58'dx;
	_BitwiseIntConcat_upper = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial _BitwiseIntConcat_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_lower = 6'dx;
	_BitwiseIntConcat_lower = 1'd0;
end
always_comb begin // combinatorial next_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_arlen = 6'dx;
	if(_chunks_are_left_D0) if(__23_D0) next_arlen = __26_D0;
	if(_chunks_are_left_D0) if(!__23_D0) next_arlen = _max_chunks_in_this_burst_D0;
end
always_comb begin // combinatorial next_last_burst_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_last_burst_in_flight = 1'bx;
	next_last_burst_in_flight = 1'b0;
	if(chunks_are_left) if(_23) next_last_burst_in_flight = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	next_last_burst_in_flight = next_last_burst_in_flight;
end
always_comb begin // combinatorial cur_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_burst_addr = 52'dx;
	cur_burst_addr = _BitwiseIntSplit_upper;
end
always_comb begin // combinatorial cur_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_align = 6'dx;
	cur_align = _BitwiseIntSplit_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_v = 58'dx;
	_BitwiseIntSplit_v = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial chunks_are_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunks_are_left = 1'bx;
	chunks_are_left = __14_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunks_are_left = chunks_are_left;
end
always_comb begin // combinatorial max_chunks_in_this_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	max_chunks_in_this_burst = 6'dx;
	if(chunks_are_left) max_chunks_in_this_burst = _18;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 33'dx;
	if(chunks_are_left) if(_23) _IntNarrow_in = __num_chunks_left_old_N1;
end
always_comb begin // combinatorial may_next_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_next_arvalid = 1'bx;
	may_next_arvalid = _39;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_next_arvalid = may_next_arvalid;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial next_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_burst_addr = 53'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) next_burst_addr = __45_D1;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_upper = 53'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_upper = next_burst_addr;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_lower = 6'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_lower = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_2_in = 59'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _IntNarrow_2_in = _BitwiseIntConcat_2_v;
end
always_comb begin // combinatorial _cur_start_chunk_addr_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_update = 1'bx;
	_cur_start_chunk_addr_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _cur_start_chunk_addr_update = 1'b1;
	if(request_new_burst) _cur_start_chunk_addr_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_update = _cur_start_chunk_addr_update;
end
always_comb begin // combinatorial _cur_start_chunk_addr_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_new = 58'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _cur_start_chunk_addr_new = _IntNarrow_2_out;
	if(_request_new_burst_D1) _cur_start_chunk_addr_new = _chunk_addr_D1;
end
always_comb begin // combinatorial next_num_chunks_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_num_chunks_left = 33'dx;
	if(!arvalid) if(may_next_arvalid) next_num_chunks_left = _IntNarrow_3_out;
end
always_comb begin // combinatorial _IntNarrow_3_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_3_in = 34'sdx;
	if(!arvalid) if(may_next_arvalid) _IntNarrow_3_in = _54;
end
always_comb begin // combinatorial _num_chunks_left_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_update = 1'bx;
	_num_chunks_left_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_update = 1'b1;
	if(request_new_burst) _num_chunks_left_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_update = _num_chunks_left_update;
end
always_comb begin // combinatorial _num_chunks_left_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_new = 33'dx;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_new = next_num_chunks_left;
	if(request_new_burst) _num_chunks_left_new = num_chunks;
end
always_comb begin // combinatorial _BoolToInt_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_i = 1'bx;
	_BoolToInt_i = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_i = _BoolToInt_i;
end
always_comb begin // combinatorial _Ternary_cond
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_cond = 1'bx;
	_Ternary_cond = _68;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Ternary_cond = _Ternary_cond;
end
always_comb begin // combinatorial _Ternary_a
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_a = 7'dx;
	_Ternary_a = _71;
end
always_comb begin // combinatorial _Ternary_b
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_b = 7'dx;
	_Ternary_b = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_4_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_4_in = 13'sdx;
	_IntNarrow_4_in = _73;
end
always_ff @(posedge aclk) begin // state final_chunk_align
	if(request_new_burst) final_chunk_align <= _BitwiseIntConcat_3_v;
end
always_ff @(posedge aclk) begin // state cur_chunk_align
	if(rvalid) cur_chunk_align <= 1'd0;
	if(request_new_burst) cur_chunk_align <= element_in_chunk_align;
end
always_comb begin // combinatorial elements_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_2 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	if(rvalid) elements_2[0] = _75;
	if(rvalid) elements_2[1] = _76;
	if(rvalid) elements_2[2] = _77;
	if(rvalid) elements_2[3] = _78;
	if(rvalid) elements_2[4] = _79;
	if(rvalid) elements_2[5] = _80;
	if(rvalid) elements_2[6] = _81;
	if(rvalid) elements_2[7] = _82;
	if(rvalid) elements_2[8] = _83;
	if(rvalid) elements_2[9] = _84;
	if(rvalid) elements_2[10] = _85;
	if(rvalid) elements_2[11] = _86;
	if(rvalid) elements_2[12] = _87;
	if(rvalid) elements_2[13] = _88;
	if(rvalid) elements_2[14] = _89;
	if(rvalid) elements_2[15] = _90;
end
always_comb begin // combinatorial num_chunk_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunk_elements = 5'dx;
	if(rvalid) if(is_last) num_chunk_elements = _IntNarrow_5_out;
	if(rvalid) if(!is_last) num_chunk_elements = _101;
end
always_comb begin // combinatorial is_last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_last = 1'bx;
	if(rvalid) is_last = _95;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_last = is_last;
end
always_comb begin // combinatorial _IntNarrow_5_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_5_in = 6'sdx;
	if(rvalid) if(is_last) _IntNarrow_5_in = _99;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _113;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial chunk_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_addr = 58'dx;
	if(request_new_burst) chunk_addr = _BitwiseIntSplit_2_upper;
end
always_comb begin // combinatorial element_in_chunk_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_in_chunk_align = 4'dx;
	if(request_new_burst) element_in_chunk_align = _BitwiseIntSplit_2_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_2_v = 62'dx;
	if(request_new_burst) _BitwiseIntSplit_2_v = _115;
end
always_comb begin // combinatorial chunk_count_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_count_bits = 33'dx;
	if(request_new_burst) chunk_count_bits = _BitwiseIntSplit_3_upper;
end
always_comb begin // combinatorial final_alignment
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	final_alignment = 4'dx;
	if(request_new_burst) final_alignment = _BitwiseIntSplit_3_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_3_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_3_v = 37'dx;
	if(request_new_burst) _BitwiseIntSplit_3_v = _118;
end
always_comb begin // combinatorial num_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunks = 33'dx;
	if(request_new_burst) if(is_no_chunks) num_chunks = 1'd1;
	if(request_new_burst) if(!is_no_chunks) num_chunks = _128;
end
always_comb begin // combinatorial is_no_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_no_chunks = 1'bx;
	if(request_new_burst) is_no_chunks = _121;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_no_chunks = is_no_chunks;
end
always_comb begin // combinatorial _BoolToInt_2_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_2_i = 1'bx;
	if(request_new_burst) if(!is_no_chunks) _BoolToInt_2_i = _127;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_2_i = _BoolToInt_2_i;
end
always_comb begin // combinatorial _BoolToInt_3_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_3_i = 1'bx;
	if(request_new_burst) _BoolToInt_3_i = _138;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_3_i = _BoolToInt_3_i;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_upper = 1'dx;
	if(request_new_burst) _BitwiseIntConcat_3_upper = _BoolToInt_3_o;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BitwiseIntConcat_3_upper = _BitwiseIntConcat_3_upper;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_lower = 4'dx;
	if(request_new_burst) _BitwiseIntConcat_3_lower = final_alignment;
end
always_comb begin // combinatorial _cur_start_chunk_addr_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_rst = 1'bx;
	_cur_start_chunk_addr_rst = _142;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_rst = _cur_start_chunk_addr_rst;
end
always_comb begin // combinatorial _num_chunks_left_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_rst = 1'bx;
	_num_chunks_left_rst = _144;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_rst = _num_chunks_left_rst;
end
endmodule

// BitwiseIntSplit #(TO: 68719476751, LOWER_BITS: 4)
module BitwiseIntSplit_TO_68719476751_LOWER_BITS_4(
	input clk,
	input wire[36:0] v,
	output /*mux_wire*/ logic[32:0] upper,
	output /*mux_wire*/ logic[3:0] lower
);

genvar _g0;
/*mux_wire*/ logic[36:0] v_bits;
/*mux_wire*/ logic[36:0] _UIntToBits_value;
wire[36:0] _UIntToBits_bits;
wire[3:0] _2;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_bits;
wire[3:0] _BitsToUInt_value;
wire[32:0] _3;
generate
for(_g0 = 0; _g0 < 33; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[4 + _g0];
end
endgenerate
/*mux_wire*/ logic[32:0] _FromBits_bits;
wire[32:0] _FromBits_value;
UIntToBits_NUM_BITS_37 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_4 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_4294967297 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 33'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 4'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 37'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 37'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 4'bxxxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// UIntToBits #(NUM_BITS: 37)
module UIntToBits_NUM_BITS_37(
	input clk,
	input wire[36:0] value,
	output /*mux_wire*/ logic[36:0] bits
);

	assign bits = value;
endmodule

// IntNarrow #(FROM_I: -64, TO_I: 4294967298, FROM: 0, TO: 4294967299)
module IntNarrow_FROM_I_64_TO_I_4294967298_FROM_0_TO_4294967299(
	input clk,
	input wire signed[33:0] in,
	output /*mux_wire*/ logic[32:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 4294967299, FROM: 1, TO: 65)
module IntNarrow_FROM_I_0_TO_I_4294967299_FROM_1_TO_65(
	input clk,
	input wire[32:0] in,
	output /*mux_wire*/ logic[6:0] out
);

	assign out = in;
endmodule

// benchmark_burst_read #(AXI_WIDTH: 256)
module benchmark_burst_read_AXI_WIDTH_256(
	input aclk,
	input wire aresetn,
	input wire[11:0] s_axi_control_awaddr,
	input wire s_axi_control_awvalid,
	output /*mux_wire*/ logic s_axi_control_awready,
	input wire[31:0] s_axi_control_wdata,
	input wire[3:0] s_axi_control_wstrb,
	input wire s_axi_control_wvalid,
	output /*mux_wire*/ logic s_axi_control_wready,
	output /*mux_wire*/ logic[1:0] s_axi_control_bresp,
	output /*mux_wire*/ logic s_axi_control_bvalid,
	input wire s_axi_control_bready,
	input wire[11:0] s_axi_control_araddr,
	input wire s_axi_control_arvalid,
	output /*mux_wire*/ logic s_axi_control_arready,
	output /*mux_wire*/ logic[31:0] s_axi_control_rdata,
	output /*mux_wire*/ logic[1:0] s_axi_control_rresp,
	output /*mux_wire*/ logic s_axi_control_rvalid,
	input wire s_axi_control_rready,
	output /*mux_wire*/ logic m_axi_awvalid,
	input wire m_axi_awready,
	output /*mux_wire*/ logic[63:0] m_axi_awaddr,
	output /*mux_wire*/ logic[7:0] m_axi_awlen,
	output /*mux_wire*/ logic[1:0] m_axi_awburst,
	output /*mux_wire*/ logic[3:0] m_axi_awcache,
	output /*mux_wire*/ logic m_axi_wvalid,
	input wire m_axi_wready,
	output /*mux_wire*/ logic[255:0] m_axi_wdata,
	output /*mux_wire*/ logic[31:0] m_axi_wstrb,
	output /*mux_wire*/ logic m_axi_wlast,
	input wire m_axi_bvalid,
	output /*mux_wire*/ logic m_axi_bready,
	input wire[1:0] m_axi_bresp,
	output /*mux_wire*/ logic m_axi_arvalid,
	input wire m_axi_arready,
	output /*mux_wire*/ logic[63:0] m_axi_araddr,
	output /*mux_wire*/ logic[7:0] m_axi_arlen,
	output /*mux_wire*/ logic[2:0] m_axi_arsize,
	output /*mux_wire*/ logic[1:0] m_axi_arburst,
	input wire m_axi_rvalid,
	output /*mux_wire*/ logic m_axi_rready,
	input wire[255:0] m_axi_rdata,
	input wire[1:0] m_axi_rresp,
	input wire m_axi_rlast,
	output /*mux_wire*/ logic[2:0] m_axi_arprot,
	output /*mux_wire*/ logic[3:0] m_axi_arcache,
	output /*mux_wire*/ logic[3:0] m_axi_arqos,
	output /*mux_wire*/ logic m_axi_arlock,
	output /*mux_wire*/ logic[3:0] m_axi_arregion
);

genvar _g0;
/*mux_wire*/ logic _ctrl_aresetn;
wire _ctrl_awready;
wire _ctrl_wready;
wire[1:0] _ctrl_bresp;
wire _ctrl_bvalid;
wire _ctrl_arready;
wire[31:0] _ctrl_rdata;
wire[1:0] _ctrl_rresp;
wire _ctrl_rvalid;
/*mux_wire*/ logic[11:0] _ctrl_awaddr;
/*mux_wire*/ logic _ctrl_awvalid;
/*mux_wire*/ logic[31:0] _ctrl_wdata;
/*mux_wire*/ logic[3:0] _ctrl_wstrb;
/*mux_wire*/ logic _ctrl_wvalid;
/*mux_wire*/ logic _ctrl_bready;
/*mux_wire*/ logic[11:0] _ctrl_araddr;
/*mux_wire*/ logic _ctrl_arvalid;
/*mux_wire*/ logic _ctrl_rready;
/*mux_wire*/ logic _reader_aresetn;
/*mux_wire*/ logic _writer_aresetn;
wire _writer_awvalid;
wire[63:0] _writer_awaddr;
wire[7:0] _writer_awlen;
wire[1:0] _writer_awburst;
wire[3:0] _writer_awcache;
wire _writer_wvalid;
wire[255:0] _writer_wdata;
wire[31:0] _writer_wstrb;
wire _writer_wlast;
wire _writer_bready;
/*mux_wire*/ logic _writer_awready;
/*mux_wire*/ logic _writer_wready;
/*mux_wire*/ logic _writer_bvalid;
/*mux_wire*/ logic[1:0] _writer_bresp;
wire _reader_arvalid;
wire[63:0] _reader_araddr;
wire[7:0] _reader_arlen;
wire[2:0] _reader_arsize;
wire[1:0] _reader_arburst;
wire _reader_rready;
/*mux_wire*/ logic _reader_arready;
/*mux_wire*/ logic _reader_rvalid;
/*mux_wire*/ logic[255:0] _reader_rdata;
/*mux_wire*/ logic[1:0] _reader_rresp;
/*mux_wire*/ logic _reader_rlast;
/*mux_wire*/ logic[63:0] addr_a_bits;
wire[31:0] _ctrl_input_regs[3:0];
wire[31:0] _46 = _ctrl_input_regs[0];
wire[31:0] _47 = _ctrl_input_regs[1];
/*mux_wire*/ logic[63:0] start_addr;
/*mux_wire*/ logic[63:0] _BitsToUInt_bits;
wire[63:0] _BitsToUInt_value;
/*mux_wire*/ logic[31:0] num_to_transfer;
wire[31:0] _49 = _ctrl_input_regs[2];
/*mux_wire*/ logic[31:0] _BitsToUInt_2_bits;
wire[31:0] _BitsToUInt_2_value;
/*mux_wire*/ logic[31:0] _IntNarrow_in;
wire[31:0] _IntNarrow_out;
/*mux_wire*/ logic[31:0] config_bits;
wire[31:0] _50 = _ctrl_input_regs[3];
wire[2:0] _51;
generate
for(_g0 = 0; _g0 < 3; _g0 = _g0 + 1) begin
assign _51[_g0] = config_bits[5 + _g0];
end
endgenerate
wire[3:0] _52;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _52[_g0] = config_bits[8 + _g0];
end
endgenerate
wire[3:0] _53;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _53[_g0] = config_bits[12 + _g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_3_bits;
wire[3:0] _BitsToUInt_3_value;
wire _54 = config_bits[16];
wire[3:0] _55;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _55[_g0] = config_bits[17 + _g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_4_bits;
wire[3:0] _BitsToUInt_4_value;
wire[10:0] _56;
generate
for(_g0 = 0; _g0 < 11; _g0 = _g0 + 1) begin
assign _56[_g0] = config_bits[21 + _g0];
end
endgenerate
/*mux_wire*/ logic[10:0] _BitsToUInt_5_bits;
wire[10:0] _BitsToUInt_5_value;
/*mux_wire*/ logic[10:0] _reader_max_in_flight;
/*state*/ logic[63:0] cycles_since_reset;
wire[64:0] _59;
assign _59 = cycles_since_reset + 1'd1;
wire[63:0] _60;
assign _60 = _59; // == mod 18446744073709551616 (target is 64 bits wide)
/*mux_wire*/ logic[63:0] cycles_since_reset_bits;
/*mux_wire*/ logic[63:0] _UIntToBits_value;
wire[63:0] _UIntToBits_bits;
/*latency*/ logic[63:0] __UIntToBits_bits_D1; always_ff @(posedge aclk) begin __UIntToBits_bits_D1 <= _UIntToBits_bits; end
/*latency*/ logic[63:0] __UIntToBits_bits_D2; always_ff @(posedge aclk) begin __UIntToBits_bits_D2 <= __UIntToBits_bits_D1; end
/*latency*/ logic[63:0] __UIntToBits_bits_D3; always_ff @(posedge aclk) begin __UIntToBits_bits_D3 <= __UIntToBits_bits_D2; end
/*state*/ logic[63:0] cycles_since_reset_at_start;
/*state*/ logic running;
/*state*/ logic[31:0] num_cycles_running;
/*state*/ logic[31:0] hash;
wire _ctrl_start;
/*latency*/ logic __ctrl_start_D1; always_ff @(posedge aclk) begin __ctrl_start_D1 <= _ctrl_start; end
/*latency*/ logic __ctrl_start_D2; always_ff @(posedge aclk) begin __ctrl_start_D2 <= __ctrl_start_D1; end
/*latency*/ logic __ctrl_start_D3; always_ff @(posedge aclk) begin __ctrl_start_D3 <= __ctrl_start_D2; end
/*mux_wire*/ logic _reader_request_new_burst;
/*mux_wire*/ logic[63:0] _reader_start_addr;
/*mux_wire*/ logic[31:0] _reader_count;
localparam[31:0] _67 = 32'b00000000000000000000000000000000;
wire[32:0] _72;
assign _72 = num_cycles_running + 1'd1;
wire[31:0] _73;
assign _73 = _72; // == mod 4294967296 (target is 32 bits wide)
/*mux_wire*/ logic _reader_is_ready_to_receive_lots_of_data;
wire _reader_value_valid;
/*latency*/ logic __reader_value_valid_D1; always_ff @(posedge aclk) begin __reader_value_valid_D1 <= _reader_value_valid; end
/*latency*/ logic __reader_value_valid_D2; always_ff @(posedge aclk) begin __reader_value_valid_D2 <= __reader_value_valid_D1; end
/*latency*/ logic __reader_value_valid_D3; always_ff @(posedge aclk) begin __reader_value_valid_D3 <= __reader_value_valid_D2; end
wire[31:0] _reader_value[7:0];
wire _reader_last;
/*mux_wire*/ logic[31:0] value[7:0];
/*mux_wire*/ logic last;
/*latency*/ logic _last_D1; always_ff @(posedge aclk) begin _last_D1 <= last; end
/*latency*/ logic _last_D2; always_ff @(posedge aclk) begin _last_D2 <= _last_D1; end
/*latency*/ logic _last_D3; always_ff @(posedge aclk) begin _last_D3 <= _last_D2; end
/*mux_wire*/ logic[31:0] new_hash_contrib;
wire[7:0] _74;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _74[_g0] = value[_g0][0];
end
endgenerate
wire _75;
assign _75 = ^_74;
/*latency*/ logic __75_D1; always_ff @(posedge aclk) begin __75_D1 <= _75; end
/*latency*/ logic __75_D2; always_ff @(posedge aclk) begin __75_D2 <= __75_D1; end
wire[7:0] _76;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _76[_g0] = value[_g0][1];
end
endgenerate
wire _77;
assign _77 = ^_76;
/*latency*/ logic __77_D1; always_ff @(posedge aclk) begin __77_D1 <= _77; end
/*latency*/ logic __77_D2; always_ff @(posedge aclk) begin __77_D2 <= __77_D1; end
wire[7:0] _78;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _78[_g0] = value[_g0][2];
end
endgenerate
wire _79;
assign _79 = ^_78;
/*latency*/ logic __79_D1; always_ff @(posedge aclk) begin __79_D1 <= _79; end
/*latency*/ logic __79_D2; always_ff @(posedge aclk) begin __79_D2 <= __79_D1; end
wire[7:0] _80;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _80[_g0] = value[_g0][3];
end
endgenerate
wire _81;
assign _81 = ^_80;
/*latency*/ logic __81_D1; always_ff @(posedge aclk) begin __81_D1 <= _81; end
/*latency*/ logic __81_D2; always_ff @(posedge aclk) begin __81_D2 <= __81_D1; end
wire[7:0] _82;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _82[_g0] = value[_g0][4];
end
endgenerate
wire _83;
assign _83 = ^_82;
/*latency*/ logic __83_D1; always_ff @(posedge aclk) begin __83_D1 <= _83; end
/*latency*/ logic __83_D2; always_ff @(posedge aclk) begin __83_D2 <= __83_D1; end
wire[7:0] _84;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _84[_g0] = value[_g0][5];
end
endgenerate
wire _85;
assign _85 = ^_84;
/*latency*/ logic __85_D1; always_ff @(posedge aclk) begin __85_D1 <= _85; end
/*latency*/ logic __85_D2; always_ff @(posedge aclk) begin __85_D2 <= __85_D1; end
wire[7:0] _86;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _86[_g0] = value[_g0][6];
end
endgenerate
wire _87;
assign _87 = ^_86;
/*latency*/ logic __87_D1; always_ff @(posedge aclk) begin __87_D1 <= _87; end
/*latency*/ logic __87_D2; always_ff @(posedge aclk) begin __87_D2 <= __87_D1; end
wire[7:0] _88;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _88[_g0] = value[_g0][7];
end
endgenerate
wire _89;
assign _89 = ^_88;
/*latency*/ logic __89_D1; always_ff @(posedge aclk) begin __89_D1 <= _89; end
/*latency*/ logic __89_D2; always_ff @(posedge aclk) begin __89_D2 <= __89_D1; end
wire[7:0] _90;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _90[_g0] = value[_g0][8];
end
endgenerate
wire _91;
assign _91 = ^_90;
/*latency*/ logic __91_D1; always_ff @(posedge aclk) begin __91_D1 <= _91; end
/*latency*/ logic __91_D2; always_ff @(posedge aclk) begin __91_D2 <= __91_D1; end
wire[7:0] _92;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _92[_g0] = value[_g0][9];
end
endgenerate
wire _93;
assign _93 = ^_92;
/*latency*/ logic __93_D1; always_ff @(posedge aclk) begin __93_D1 <= _93; end
/*latency*/ logic __93_D2; always_ff @(posedge aclk) begin __93_D2 <= __93_D1; end
wire[7:0] _94;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _94[_g0] = value[_g0][10];
end
endgenerate
wire _95;
assign _95 = ^_94;
/*latency*/ logic __95_D1; always_ff @(posedge aclk) begin __95_D1 <= _95; end
/*latency*/ logic __95_D2; always_ff @(posedge aclk) begin __95_D2 <= __95_D1; end
wire[7:0] _96;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _96[_g0] = value[_g0][11];
end
endgenerate
wire _97;
assign _97 = ^_96;
/*latency*/ logic __97_D1; always_ff @(posedge aclk) begin __97_D1 <= _97; end
/*latency*/ logic __97_D2; always_ff @(posedge aclk) begin __97_D2 <= __97_D1; end
wire[7:0] _98;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _98[_g0] = value[_g0][12];
end
endgenerate
wire _99;
assign _99 = ^_98;
/*latency*/ logic __99_D1; always_ff @(posedge aclk) begin __99_D1 <= _99; end
/*latency*/ logic __99_D2; always_ff @(posedge aclk) begin __99_D2 <= __99_D1; end
wire[7:0] _100;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _100[_g0] = value[_g0][13];
end
endgenerate
wire _101;
assign _101 = ^_100;
/*latency*/ logic __101_D1; always_ff @(posedge aclk) begin __101_D1 <= _101; end
/*latency*/ logic __101_D2; always_ff @(posedge aclk) begin __101_D2 <= __101_D1; end
wire[7:0] _102;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _102[_g0] = value[_g0][14];
end
endgenerate
wire _103;
assign _103 = ^_102;
/*latency*/ logic __103_D1; always_ff @(posedge aclk) begin __103_D1 <= _103; end
/*latency*/ logic __103_D2; always_ff @(posedge aclk) begin __103_D2 <= __103_D1; end
wire[7:0] _104;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _104[_g0] = value[_g0][15];
end
endgenerate
wire _105;
assign _105 = ^_104;
/*latency*/ logic __105_D1; always_ff @(posedge aclk) begin __105_D1 <= _105; end
/*latency*/ logic __105_D2; always_ff @(posedge aclk) begin __105_D2 <= __105_D1; end
wire[7:0] _106;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _106[_g0] = value[_g0][16];
end
endgenerate
wire _107;
assign _107 = ^_106;
/*latency*/ logic __107_D1; always_ff @(posedge aclk) begin __107_D1 <= _107; end
/*latency*/ logic __107_D2; always_ff @(posedge aclk) begin __107_D2 <= __107_D1; end
wire[7:0] _108;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _108[_g0] = value[_g0][17];
end
endgenerate
wire _109;
assign _109 = ^_108;
/*latency*/ logic __109_D1; always_ff @(posedge aclk) begin __109_D1 <= _109; end
/*latency*/ logic __109_D2; always_ff @(posedge aclk) begin __109_D2 <= __109_D1; end
wire[7:0] _110;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _110[_g0] = value[_g0][18];
end
endgenerate
wire _111;
assign _111 = ^_110;
/*latency*/ logic __111_D1; always_ff @(posedge aclk) begin __111_D1 <= _111; end
/*latency*/ logic __111_D2; always_ff @(posedge aclk) begin __111_D2 <= __111_D1; end
wire[7:0] _112;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _112[_g0] = value[_g0][19];
end
endgenerate
wire _113;
assign _113 = ^_112;
/*latency*/ logic __113_D1; always_ff @(posedge aclk) begin __113_D1 <= _113; end
/*latency*/ logic __113_D2; always_ff @(posedge aclk) begin __113_D2 <= __113_D1; end
wire[7:0] _114;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _114[_g0] = value[_g0][20];
end
endgenerate
wire _115;
assign _115 = ^_114;
/*latency*/ logic __115_D1; always_ff @(posedge aclk) begin __115_D1 <= _115; end
/*latency*/ logic __115_D2; always_ff @(posedge aclk) begin __115_D2 <= __115_D1; end
wire[7:0] _116;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _116[_g0] = value[_g0][21];
end
endgenerate
wire _117;
assign _117 = ^_116;
/*latency*/ logic __117_D1; always_ff @(posedge aclk) begin __117_D1 <= _117; end
/*latency*/ logic __117_D2; always_ff @(posedge aclk) begin __117_D2 <= __117_D1; end
wire[7:0] _118;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _118[_g0] = value[_g0][22];
end
endgenerate
wire _119;
assign _119 = ^_118;
/*latency*/ logic __119_D1; always_ff @(posedge aclk) begin __119_D1 <= _119; end
/*latency*/ logic __119_D2; always_ff @(posedge aclk) begin __119_D2 <= __119_D1; end
wire[7:0] _120;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _120[_g0] = value[_g0][23];
end
endgenerate
wire _121;
assign _121 = ^_120;
/*latency*/ logic __121_D1; always_ff @(posedge aclk) begin __121_D1 <= _121; end
/*latency*/ logic __121_D2; always_ff @(posedge aclk) begin __121_D2 <= __121_D1; end
wire[7:0] _122;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _122[_g0] = value[_g0][24];
end
endgenerate
wire _123;
assign _123 = ^_122;
/*latency*/ logic __123_D1; always_ff @(posedge aclk) begin __123_D1 <= _123; end
/*latency*/ logic __123_D2; always_ff @(posedge aclk) begin __123_D2 <= __123_D1; end
wire[7:0] _124;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _124[_g0] = value[_g0][25];
end
endgenerate
wire _125;
assign _125 = ^_124;
/*latency*/ logic __125_D1; always_ff @(posedge aclk) begin __125_D1 <= _125; end
/*latency*/ logic __125_D2; always_ff @(posedge aclk) begin __125_D2 <= __125_D1; end
wire[7:0] _126;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _126[_g0] = value[_g0][26];
end
endgenerate
wire _127;
assign _127 = ^_126;
/*latency*/ logic __127_D1; always_ff @(posedge aclk) begin __127_D1 <= _127; end
/*latency*/ logic __127_D2; always_ff @(posedge aclk) begin __127_D2 <= __127_D1; end
wire[7:0] _128;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _128[_g0] = value[_g0][27];
end
endgenerate
wire _129;
assign _129 = ^_128;
/*latency*/ logic __129_D1; always_ff @(posedge aclk) begin __129_D1 <= _129; end
/*latency*/ logic __129_D2; always_ff @(posedge aclk) begin __129_D2 <= __129_D1; end
wire[7:0] _130;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _130[_g0] = value[_g0][28];
end
endgenerate
wire _131;
assign _131 = ^_130;
/*latency*/ logic __131_D1; always_ff @(posedge aclk) begin __131_D1 <= _131; end
/*latency*/ logic __131_D2; always_ff @(posedge aclk) begin __131_D2 <= __131_D1; end
wire[7:0] _132;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _132[_g0] = value[_g0][29];
end
endgenerate
wire _133;
assign _133 = ^_132;
/*latency*/ logic __133_D1; always_ff @(posedge aclk) begin __133_D1 <= _133; end
/*latency*/ logic __133_D2; always_ff @(posedge aclk) begin __133_D2 <= __133_D1; end
wire[7:0] _134;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _134[_g0] = value[_g0][30];
end
endgenerate
wire _135;
assign _135 = ^_134;
/*latency*/ logic __135_D1; always_ff @(posedge aclk) begin __135_D1 <= _135; end
/*latency*/ logic __135_D2; always_ff @(posedge aclk) begin __135_D2 <= __135_D1; end
wire[7:0] _136;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _136[_g0] = value[_g0][31];
end
endgenerate
wire _137;
assign _137 = ^_136;
/*latency*/ logic __137_D1; always_ff @(posedge aclk) begin __137_D1 <= _137; end
/*latency*/ logic __137_D2; always_ff @(posedge aclk) begin __137_D2 <= __137_D1; end
/*mux_wire*/ logic[31:0] new_hash;
/*latency*/ logic[31:0] _new_hash_D3; always_ff @(posedge aclk) begin _new_hash_D3 <= new_hash; end
wire[31:0] _140;
assign _140 = hash ^ new_hash_contrib;
/*mux_wire*/ logic[31:0] _UIntToBits_2_value;
wire[31:0] _UIntToBits_2_bits;
/*latency*/ logic[31:0] __UIntToBits_2_bits_D1; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D1 <= _UIntToBits_2_bits; end
/*latency*/ logic[31:0] __UIntToBits_2_bits_D2; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D2 <= __UIntToBits_2_bits_D1; end
/*latency*/ logic[31:0] __UIntToBits_2_bits_D3; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D3 <= __UIntToBits_2_bits_D2; end
wire[31:0] _144;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _144[_g0] = cycles_since_reset_at_start[_g0];
end
endgenerate
wire[31:0] _145;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _145[_g0] = cycles_since_reset_at_start[32 + _g0];
end
endgenerate
wire[31:0] _146;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _146[_g0] = cycles_since_reset_bits[_g0];
end
endgenerate
wire[31:0] _147;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _147[_g0] = cycles_since_reset_bits[32 + _g0];
end
endgenerate
wire[31:0] _148[5:0];
assign _148[0] = __UIntToBits_2_bits_D3;
assign _148[1] = _new_hash_D3;
assign _148[2] = _144;
assign _148[3] = _145;
assign _148[4] = _146;
assign _148[5] = _147;
/*mux_wire*/ logic _ctrl_finish;
/*mux_wire*/ logic[31:0] _ctrl_output_regs[5:0];
wire _153;
assign _153 = !aresetn;
/*latency*/ logic __153_D1; always_ff @(posedge aclk) begin __153_D1 <= _153; end
/*latency*/ logic __153_D2; always_ff @(posedge aclk) begin __153_D2 <= __153_D1; end
localparam[31:0] _155 = 32'b00000000000000000000000000000000;
axi_ctrl_slave_NUM_INPUT_REGS_4_NUM_OUTPUT_REGS_6_ADDR_WIDTH_12_AXI_WIDTH_32 ctrl(
	.aclk(aclk),
	.aresetn(_ctrl_aresetn),
	.awaddr(_ctrl_awaddr),
	.awvalid(_ctrl_awvalid),
	.awready(_ctrl_awready),
	.wdata(_ctrl_wdata),
	.wstrb(_ctrl_wstrb),
	.wvalid(_ctrl_wvalid),
	.wready(_ctrl_wready),
	.bresp(_ctrl_bresp),
	.bvalid(_ctrl_bvalid),
	.bready(_ctrl_bready),
	.araddr(_ctrl_araddr),
	.arvalid(_ctrl_arvalid),
	.arready(_ctrl_arready),
	.rdata(_ctrl_rdata),
	.rresp(_ctrl_rresp),
	.rvalid(_ctrl_rvalid),
	.rready(_ctrl_rready),
	.input_regs(_ctrl_input_regs),
	.start(_ctrl_start),
	.finish(_ctrl_finish),
	.output_regs(_ctrl_output_regs)
);
axi_realigning_burst_reader_T_type_bool_32_8_AXI_WIDTH_256_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616 reader(
	.aclk(aclk),
	.aresetn(_reader_aresetn),
	.arvalid(_reader_arvalid),
	.arready(_reader_arready),
	.araddr(_reader_araddr),
	.arlen(_reader_arlen),
	.arsize(_reader_arsize),
	.arburst(_reader_arburst),
	.arprot(),
	.arcache(),
	.arqos(),
	.arlock(),
	.arregion(),
	.rvalid(_reader_rvalid),
	.rready(_reader_rready),
	.rdata(_reader_rdata),
	.rresp(_reader_rresp),
	.rlast(_reader_rlast),
	.max_in_flight(_reader_max_in_flight),
	.may_request_new_burst(),
	.request_new_burst(_reader_request_new_burst),
	.start_addr(_reader_start_addr),
	.count(_reader_count),
	.is_ready_to_receive_lots_of_data(_reader_is_ready_to_receive_lots_of_data),
	.value_valid(_reader_value_valid),
	.value(_reader_value),
	.last(_reader_last)
);
axi_memory_writer_tie_off_AXI_WIDTH_256 writer(
	.aclk(aclk),
	.aresetn(_writer_aresetn),
	.awvalid(_writer_awvalid),
	.awready(_writer_awready),
	.awaddr(_writer_awaddr),
	.awlen(_writer_awlen),
	.awsize(),
	.awburst(_writer_awburst),
	.awprot(),
	.awcache(_writer_awcache),
	.awqos(),
	.awlock(),
	.awregion(),
	.wvalid(_writer_wvalid),
	.wready(_writer_wready),
	.wdata(_writer_wdata),
	.wstrb(_writer_wstrb),
	.wlast(_writer_wlast),
	.bvalid(_writer_bvalid),
	.bresp(_writer_bresp),
	.bready(_writer_bready)
);
BitsToUInt_NUM_BITS_64 BitsToUInt(
	.clk(aclk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
BitsToUInt_NUM_BITS_32 BitsToUInt_2(
	.clk(aclk),
	.bits(_BitsToUInt_2_bits),
	.value(_BitsToUInt_2_value)
);
IntNarrow_FROM_I_0_TO_I_4294967296_FROM_1_TO_4294967296 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
BitsToUInt_NUM_BITS_4 BitsToUInt_3(
	.clk(aclk),
	.bits(_BitsToUInt_3_bits),
	.value(_BitsToUInt_3_value)
);
BitsToUInt_NUM_BITS_4 BitsToUInt_4(
	.clk(aclk),
	.bits(_BitsToUInt_4_bits),
	.value(_BitsToUInt_4_value)
);
BitsToUInt_NUM_BITS_11 BitsToUInt_5(
	.clk(aclk),
	.bits(_BitsToUInt_5_bits),
	.value(_BitsToUInt_5_value)
);
UIntToBits_NUM_BITS_64 UIntToBits(
	.clk(aclk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_32 UIntToBits_2(
	.clk(aclk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
always_comb begin // combinatorial _ctrl_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_aresetn = 1'bx;
	_ctrl_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_aresetn = _ctrl_aresetn;
end
always_comb begin // combinatorial s_axi_control_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_awready = 1'bx;
	s_axi_control_awready = _ctrl_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_awready = s_axi_control_awready;
end
always_comb begin // combinatorial s_axi_control_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_wready = 1'bx;
	s_axi_control_wready = _ctrl_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_wready = s_axi_control_wready;
end
always_comb begin // combinatorial s_axi_control_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bresp = 2'bxx;
	s_axi_control_bresp = _ctrl_bresp;
end
always_comb begin // combinatorial s_axi_control_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bvalid = 1'bx;
	s_axi_control_bvalid = _ctrl_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_bvalid = s_axi_control_bvalid;
end
always_comb begin // combinatorial s_axi_control_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_arready = 1'bx;
	s_axi_control_arready = _ctrl_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_arready = s_axi_control_arready;
end
always_comb begin // combinatorial s_axi_control_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	s_axi_control_rdata = _ctrl_rdata;
end
always_comb begin // combinatorial s_axi_control_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rresp = 2'bxx;
	s_axi_control_rresp = _ctrl_rresp;
end
always_comb begin // combinatorial s_axi_control_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rvalid = 1'bx;
	s_axi_control_rvalid = _ctrl_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_rvalid = s_axi_control_rvalid;
end
always_comb begin // combinatorial _ctrl_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awaddr = 12'dx;
	_ctrl_awaddr = s_axi_control_awaddr;
end
always_comb begin // combinatorial _ctrl_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awvalid = 1'bx;
	_ctrl_awvalid = s_axi_control_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_awvalid = _ctrl_awvalid;
end
always_comb begin // combinatorial _ctrl_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_ctrl_wdata = s_axi_control_wdata;
end
always_comb begin // combinatorial _ctrl_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wstrb = 4'bxxxx;
	_ctrl_wstrb = s_axi_control_wstrb;
end
always_comb begin // combinatorial _ctrl_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wvalid = 1'bx;
	_ctrl_wvalid = s_axi_control_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_wvalid = _ctrl_wvalid;
end
always_comb begin // combinatorial _ctrl_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_bready = 1'bx;
	_ctrl_bready = s_axi_control_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_bready = _ctrl_bready;
end
always_comb begin // combinatorial _ctrl_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_araddr = 12'dx;
	_ctrl_araddr = s_axi_control_araddr;
end
always_comb begin // combinatorial _ctrl_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_arvalid = 1'bx;
	_ctrl_arvalid = s_axi_control_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_arvalid = _ctrl_arvalid;
end
always_comb begin // combinatorial _ctrl_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_rready = 1'bx;
	_ctrl_rready = s_axi_control_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_rready = _ctrl_rready;
end
always_comb begin // combinatorial _reader_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_aresetn = 1'bx;
	_reader_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_aresetn = _reader_aresetn;
end
always_comb begin // combinatorial _writer_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_aresetn = 1'bx;
	_writer_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_aresetn = _writer_aresetn;
end
always_comb begin // combinatorial m_axi_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awvalid = 1'bx;
	m_axi_awvalid = _writer_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_awvalid = m_axi_awvalid;
end
always_comb begin // combinatorial m_axi_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awaddr = 64'dx;
	m_axi_awaddr = _writer_awaddr;
end
always_comb begin // combinatorial m_axi_awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awlen = 8'dx;
	m_axi_awlen = _writer_awlen;
end
always_comb begin // combinatorial m_axi_awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awburst = 2'bxx;
	m_axi_awburst = _writer_awburst;
end
always_comb begin // combinatorial m_axi_awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awcache = 4'bxxxx;
	m_axi_awcache = _writer_awcache;
end
always_comb begin // combinatorial m_axi_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wvalid = 1'bx;
	m_axi_wvalid = _writer_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wvalid = m_axi_wvalid;
end
always_comb begin // combinatorial m_axi_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wdata = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	m_axi_wdata = _writer_wdata;
end
always_comb begin // combinatorial m_axi_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wstrb = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	m_axi_wstrb = _writer_wstrb;
end
always_comb begin // combinatorial m_axi_wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wlast = 1'bx;
	m_axi_wlast = _writer_wlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wlast = m_axi_wlast;
end
always_comb begin // combinatorial m_axi_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_bready = 1'bx;
	m_axi_bready = _writer_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_bready = m_axi_bready;
end
always_comb begin // combinatorial _writer_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_awready = 1'bx;
	_writer_awready = m_axi_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_awready = _writer_awready;
end
always_comb begin // combinatorial _writer_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_wready = 1'bx;
	_writer_wready = m_axi_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_wready = _writer_wready;
end
always_comb begin // combinatorial _writer_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bvalid = 1'bx;
	_writer_bvalid = m_axi_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_bvalid = _writer_bvalid;
end
always_comb begin // combinatorial _writer_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bresp = 2'bxx;
	_writer_bresp = m_axi_bresp;
end
always_comb begin // combinatorial m_axi_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arvalid = 1'bx;
	m_axi_arvalid = _reader_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arvalid = m_axi_arvalid;
end
always_comb begin // combinatorial m_axi_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_araddr = 64'dx;
	m_axi_araddr = _reader_araddr;
end
always_comb begin // combinatorial m_axi_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlen = 8'dx;
	m_axi_arlen = _reader_arlen;
end
always_comb begin // combinatorial m_axi_arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arsize = 3'dx;
	m_axi_arsize = _reader_arsize;
end
always_comb begin // combinatorial m_axi_arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arburst = 2'bxx;
	m_axi_arburst = _reader_arburst;
end
always_comb begin // combinatorial m_axi_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_rready = 1'bx;
	m_axi_rready = _reader_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_rready = m_axi_rready;
end
always_comb begin // combinatorial _reader_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_arready = 1'bx;
	_reader_arready = m_axi_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_arready = _reader_arready;
end
always_comb begin // combinatorial _reader_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rvalid = 1'bx;
	_reader_rvalid = m_axi_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rvalid = _reader_rvalid;
end
always_comb begin // combinatorial _reader_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rdata = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_reader_rdata = m_axi_rdata;
end
always_comb begin // combinatorial _reader_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rresp = 2'bxx;
	_reader_rresp = m_axi_rresp;
end
always_comb begin // combinatorial _reader_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rlast = 1'bx;
	_reader_rlast = m_axi_rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rlast = _reader_rlast;
end
always_comb begin // combinatorial addr_a_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	addr_a_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[_v0] = _46[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[32 + _v0] = _47[_v0];
end
end
always_comb begin // combinatorial start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	start_addr = 64'dx;
	start_addr = _BitsToUInt_value;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_BitsToUInt_bits = addr_a_bits;
end
always_comb begin // combinatorial num_to_transfer
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_to_transfer = 32'dx;
	num_to_transfer = _IntNarrow_out;
end
always_comb begin // combinatorial _BitsToUInt_2_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_2_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_BitsToUInt_2_bits = _49;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 32'dx;
	_IntNarrow_in = _BitsToUInt_2_value;
end
always_comb begin // combinatorial config_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	config_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	config_bits = _50;
end
always_comb begin // combinatorial m_axi_arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arprot = 3'bxxx;
	m_axi_arprot = _51;
end
always_comb begin // combinatorial m_axi_arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arcache = 4'bxxxx;
	m_axi_arcache = _52;
end
always_comb begin // combinatorial m_axi_arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arqos = 4'dx;
	m_axi_arqos = _BitsToUInt_3_value;
end
always_comb begin // combinatorial _BitsToUInt_3_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_3_bits = 4'bxxxx;
	_BitsToUInt_3_bits = _53;
end
always_comb begin // combinatorial m_axi_arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlock = 1'bx;
	m_axi_arlock = _54;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arlock = m_axi_arlock;
end
always_comb begin // combinatorial m_axi_arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arregion = 4'dx;
	m_axi_arregion = _BitsToUInt_4_value;
end
always_comb begin // combinatorial _BitsToUInt_4_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_4_bits = 4'bxxxx;
	_BitsToUInt_4_bits = _55;
end
always_comb begin // combinatorial _BitsToUInt_5_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_5_bits = 11'bxxxxxxxxxxx;
	_BitsToUInt_5_bits = _56;
end
always_comb begin // combinatorial _reader_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_max_in_flight = 11'dx;
	_reader_max_in_flight = _BitsToUInt_5_value;
end
always_ff @(posedge aclk) begin // state cycles_since_reset
	cycles_since_reset <= _60;
	if(_153) cycles_since_reset <= 1'd0;
end
always_comb begin // combinatorial cycles_since_reset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cycles_since_reset_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	cycles_since_reset_bits = __UIntToBits_bits_D3;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 64'dx;
	_UIntToBits_value = cycles_since_reset;
end
always_ff @(posedge aclk) begin // state cycles_since_reset_at_start
	if(__ctrl_start_D3) cycles_since_reset_at_start <= cycles_since_reset_bits;
end
always_ff @(posedge aclk) begin // state running
	if(_ctrl_start) running <= 1'b1;
	if(_reader_value_valid) if(last) running <= 1'b0;
	if(_153) running <= 1'b0;
end
always_ff @(posedge aclk) begin // state num_cycles_running
	if(_ctrl_start) num_cycles_running <= 1'd0;
	if(running) num_cycles_running <= _73;
	if(_153) num_cycles_running <= 1'd0;
end
always_ff @(posedge aclk) begin // state hash
	if(__ctrl_start_D2) hash <= _67;
	if(__reader_value_valid_D2) hash <= new_hash;
	if(__153_D2) hash <= _155;
end
always_comb begin // combinatorial _reader_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_request_new_burst = 1'bx;
	_reader_request_new_burst = 1'b0;
	if(_ctrl_start) _reader_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_request_new_burst = _reader_request_new_burst;
end
always_comb begin // combinatorial _reader_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_start_addr = 64'dx;
	if(_ctrl_start) _reader_start_addr = start_addr;
end
always_comb begin // combinatorial _reader_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_count = 32'dx;
	if(_ctrl_start) _reader_count = num_to_transfer;
end
always_comb begin // combinatorial _reader_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_is_ready_to_receive_lots_of_data = 1'bx;
	_reader_is_ready_to_receive_lots_of_data = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_is_ready_to_receive_lots_of_data = _reader_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_reader_value_valid) value[_v0] = _reader_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_reader_value_valid) last = _reader_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_comb begin // combinatorial new_hash_contrib
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_hash_contrib = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(__reader_value_valid_D2) new_hash_contrib[0] = __75_D2;
	if(__reader_value_valid_D2) new_hash_contrib[1] = __77_D2;
	if(__reader_value_valid_D2) new_hash_contrib[2] = __79_D2;
	if(__reader_value_valid_D2) new_hash_contrib[3] = __81_D2;
	if(__reader_value_valid_D2) new_hash_contrib[4] = __83_D2;
	if(__reader_value_valid_D2) new_hash_contrib[5] = __85_D2;
	if(__reader_value_valid_D2) new_hash_contrib[6] = __87_D2;
	if(__reader_value_valid_D2) new_hash_contrib[7] = __89_D2;
	if(__reader_value_valid_D2) new_hash_contrib[8] = __91_D2;
	if(__reader_value_valid_D2) new_hash_contrib[9] = __93_D2;
	if(__reader_value_valid_D2) new_hash_contrib[10] = __95_D2;
	if(__reader_value_valid_D2) new_hash_contrib[11] = __97_D2;
	if(__reader_value_valid_D2) new_hash_contrib[12] = __99_D2;
	if(__reader_value_valid_D2) new_hash_contrib[13] = __101_D2;
	if(__reader_value_valid_D2) new_hash_contrib[14] = __103_D2;
	if(__reader_value_valid_D2) new_hash_contrib[15] = __105_D2;
	if(__reader_value_valid_D2) new_hash_contrib[16] = __107_D2;
	if(__reader_value_valid_D2) new_hash_contrib[17] = __109_D2;
	if(__reader_value_valid_D2) new_hash_contrib[18] = __111_D2;
	if(__reader_value_valid_D2) new_hash_contrib[19] = __113_D2;
	if(__reader_value_valid_D2) new_hash_contrib[20] = __115_D2;
	if(__reader_value_valid_D2) new_hash_contrib[21] = __117_D2;
	if(__reader_value_valid_D2) new_hash_contrib[22] = __119_D2;
	if(__reader_value_valid_D2) new_hash_contrib[23] = __121_D2;
	if(__reader_value_valid_D2) new_hash_contrib[24] = __123_D2;
	if(__reader_value_valid_D2) new_hash_contrib[25] = __125_D2;
	if(__reader_value_valid_D2) new_hash_contrib[26] = __127_D2;
	if(__reader_value_valid_D2) new_hash_contrib[27] = __129_D2;
	if(__reader_value_valid_D2) new_hash_contrib[28] = __131_D2;
	if(__reader_value_valid_D2) new_hash_contrib[29] = __133_D2;
	if(__reader_value_valid_D2) new_hash_contrib[30] = __135_D2;
	if(__reader_value_valid_D2) new_hash_contrib[31] = __137_D2;
end
always_comb begin // combinatorial new_hash
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_hash = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(__reader_value_valid_D2) new_hash = _140;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 32'dx;
	if(_reader_value_valid) if(last) _UIntToBits_2_value = num_cycles_running;
end
always_comb begin // combinatorial _ctrl_finish
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_finish = 1'bx;
	_ctrl_finish = 1'b0;
	if(__reader_value_valid_D3) if(_last_D3) _ctrl_finish = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_finish = _ctrl_finish;
end
always_comb begin // combinatorial _ctrl_output_regs
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_output_regs = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
if(__reader_value_valid_D3) if(_last_D3) _ctrl_output_regs[_v0] = _148[_v0];
end
end
endmodule

// axi_memory_writer_tie_off #(AXI_WIDTH: 256)
module axi_memory_writer_tie_off_AXI_WIDTH_256(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic awvalid,
	input wire awready,
	output /*mux_wire*/ logic[63:0] awaddr,
	output /*mux_wire*/ logic[7:0] awlen,
	output /*mux_wire*/ logic[2:0] awsize,
	output /*mux_wire*/ logic[1:0] awburst,
	output /*mux_wire*/ logic[2:0] awprot,
	output /*mux_wire*/ logic[3:0] awcache,
	output /*mux_wire*/ logic[3:0] awqos,
	output /*mux_wire*/ logic awlock,
	output /*mux_wire*/ logic[3:0] awregion,
	output /*mux_wire*/ logic wvalid,
	input wire wready,
	output /*mux_wire*/ logic[255:0] wdata,
	output /*mux_wire*/ logic[31:0] wstrb,
	output /*mux_wire*/ logic wlast,
	input wire bvalid,
	input wire[1:0] bresp,
	output /*mux_wire*/ logic bready
);

/*mux_wire*/ logic _aresetn;
localparam[1:0] _4 = 2'b00;
localparam[2:0] _5 = 3'b000;
localparam[3:0] _6 = 4'b0000;
/*mux_wire*/ logic _Repeat_v;
wire[255:0] _Repeat_result;
/*mux_wire*/ logic _Repeat_2_v;
wire[31:0] _Repeat_2_result;
/*mux_wire*/ logic _awready;
/*mux_wire*/ logic _wready;
/*mux_wire*/ logic _bvalid;
/*mux_wire*/ logic[1:0] _bresp;
Repeat_T_type_bool_SIZE_256 Repeat(
	.clk(aclk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
Repeat_T_type_bool_SIZE_32 Repeat_2(
	.clk(aclk),
	.v(_Repeat_2_v),
	.result(_Repeat_2_result)
);
always_comb begin // combinatorial _aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_aresetn = 1'bx;
	_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_aresetn = _aresetn;
end
always_comb begin // combinatorial awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awvalid = 1'bx;
	awvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awvalid = awvalid;
end
always_comb begin // combinatorial awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awaddr = 64'dx;
	awaddr = 1'd0;
end
always_comb begin // combinatorial awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlen = 8'dx;
	awlen = 1'd0;
end
always_comb begin // combinatorial awsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awsize = 3'dx;
	awsize = 3'd5;
end
always_comb begin // combinatorial awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awburst = 2'bxx;
	awburst = _4;
end
always_comb begin // combinatorial awprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awprot = 3'bxxx;
	awprot = _5;
end
always_comb begin // combinatorial awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awcache = 4'bxxxx;
	awcache = _6;
end
always_comb begin // combinatorial awqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awqos = 4'dx;
	awqos = 1'd0;
end
always_comb begin // combinatorial awlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlock = 1'bx;
	awlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awlock = awlock;
end
always_comb begin // combinatorial awregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awregion = 4'dx;
	awregion = 1'd0;
end
always_comb begin // combinatorial wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wvalid = 1'bx;
	wvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wvalid = wvalid;
end
always_comb begin // combinatorial wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wdata = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	wdata = _Repeat_result;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	_Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
always_comb begin // combinatorial wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wstrb = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	wstrb = _Repeat_2_result;
end
always_comb begin // combinatorial _Repeat_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_2_v = 1'bx;
	_Repeat_2_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_2_v = _Repeat_2_v;
end
always_comb begin // combinatorial wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wlast = 1'bx;
	wlast = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wlast = wlast;
end
always_comb begin // combinatorial bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	bready = 1'bx;
	bready = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	bready = bready;
end
always_comb begin // combinatorial _awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_awready = 1'bx;
	_awready = awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_awready = _awready;
end
always_comb begin // combinatorial _wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_wready = 1'bx;
	_wready = wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_wready = _wready;
end
always_comb begin // combinatorial _bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_bvalid = 1'bx;
	_bvalid = bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_bvalid = _bvalid;
end
always_comb begin // combinatorial _bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_bresp = 2'bxx;
	_bresp = bresp;
end
endmodule

// Repeat #(T: type bool #(), SIZE: 256)
module Repeat_T_type_bool_SIZE_256(
	input clk,
	input wire v,
	output /*mux_wire*/ logic[255:0] result
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
	result[4] = v;
	result[5] = v;
	result[6] = v;
	result[7] = v;
	result[8] = v;
	result[9] = v;
	result[10] = v;
	result[11] = v;
	result[12] = v;
	result[13] = v;
	result[14] = v;
	result[15] = v;
	result[16] = v;
	result[17] = v;
	result[18] = v;
	result[19] = v;
	result[20] = v;
	result[21] = v;
	result[22] = v;
	result[23] = v;
	result[24] = v;
	result[25] = v;
	result[26] = v;
	result[27] = v;
	result[28] = v;
	result[29] = v;
	result[30] = v;
	result[31] = v;
	result[32] = v;
	result[33] = v;
	result[34] = v;
	result[35] = v;
	result[36] = v;
	result[37] = v;
	result[38] = v;
	result[39] = v;
	result[40] = v;
	result[41] = v;
	result[42] = v;
	result[43] = v;
	result[44] = v;
	result[45] = v;
	result[46] = v;
	result[47] = v;
	result[48] = v;
	result[49] = v;
	result[50] = v;
	result[51] = v;
	result[52] = v;
	result[53] = v;
	result[54] = v;
	result[55] = v;
	result[56] = v;
	result[57] = v;
	result[58] = v;
	result[59] = v;
	result[60] = v;
	result[61] = v;
	result[62] = v;
	result[63] = v;
	result[64] = v;
	result[65] = v;
	result[66] = v;
	result[67] = v;
	result[68] = v;
	result[69] = v;
	result[70] = v;
	result[71] = v;
	result[72] = v;
	result[73] = v;
	result[74] = v;
	result[75] = v;
	result[76] = v;
	result[77] = v;
	result[78] = v;
	result[79] = v;
	result[80] = v;
	result[81] = v;
	result[82] = v;
	result[83] = v;
	result[84] = v;
	result[85] = v;
	result[86] = v;
	result[87] = v;
	result[88] = v;
	result[89] = v;
	result[90] = v;
	result[91] = v;
	result[92] = v;
	result[93] = v;
	result[94] = v;
	result[95] = v;
	result[96] = v;
	result[97] = v;
	result[98] = v;
	result[99] = v;
	result[100] = v;
	result[101] = v;
	result[102] = v;
	result[103] = v;
	result[104] = v;
	result[105] = v;
	result[106] = v;
	result[107] = v;
	result[108] = v;
	result[109] = v;
	result[110] = v;
	result[111] = v;
	result[112] = v;
	result[113] = v;
	result[114] = v;
	result[115] = v;
	result[116] = v;
	result[117] = v;
	result[118] = v;
	result[119] = v;
	result[120] = v;
	result[121] = v;
	result[122] = v;
	result[123] = v;
	result[124] = v;
	result[125] = v;
	result[126] = v;
	result[127] = v;
	result[128] = v;
	result[129] = v;
	result[130] = v;
	result[131] = v;
	result[132] = v;
	result[133] = v;
	result[134] = v;
	result[135] = v;
	result[136] = v;
	result[137] = v;
	result[138] = v;
	result[139] = v;
	result[140] = v;
	result[141] = v;
	result[142] = v;
	result[143] = v;
	result[144] = v;
	result[145] = v;
	result[146] = v;
	result[147] = v;
	result[148] = v;
	result[149] = v;
	result[150] = v;
	result[151] = v;
	result[152] = v;
	result[153] = v;
	result[154] = v;
	result[155] = v;
	result[156] = v;
	result[157] = v;
	result[158] = v;
	result[159] = v;
	result[160] = v;
	result[161] = v;
	result[162] = v;
	result[163] = v;
	result[164] = v;
	result[165] = v;
	result[166] = v;
	result[167] = v;
	result[168] = v;
	result[169] = v;
	result[170] = v;
	result[171] = v;
	result[172] = v;
	result[173] = v;
	result[174] = v;
	result[175] = v;
	result[176] = v;
	result[177] = v;
	result[178] = v;
	result[179] = v;
	result[180] = v;
	result[181] = v;
	result[182] = v;
	result[183] = v;
	result[184] = v;
	result[185] = v;
	result[186] = v;
	result[187] = v;
	result[188] = v;
	result[189] = v;
	result[190] = v;
	result[191] = v;
	result[192] = v;
	result[193] = v;
	result[194] = v;
	result[195] = v;
	result[196] = v;
	result[197] = v;
	result[198] = v;
	result[199] = v;
	result[200] = v;
	result[201] = v;
	result[202] = v;
	result[203] = v;
	result[204] = v;
	result[205] = v;
	result[206] = v;
	result[207] = v;
	result[208] = v;
	result[209] = v;
	result[210] = v;
	result[211] = v;
	result[212] = v;
	result[213] = v;
	result[214] = v;
	result[215] = v;
	result[216] = v;
	result[217] = v;
	result[218] = v;
	result[219] = v;
	result[220] = v;
	result[221] = v;
	result[222] = v;
	result[223] = v;
	result[224] = v;
	result[225] = v;
	result[226] = v;
	result[227] = v;
	result[228] = v;
	result[229] = v;
	result[230] = v;
	result[231] = v;
	result[232] = v;
	result[233] = v;
	result[234] = v;
	result[235] = v;
	result[236] = v;
	result[237] = v;
	result[238] = v;
	result[239] = v;
	result[240] = v;
	result[241] = v;
	result[242] = v;
	result[243] = v;
	result[244] = v;
	result[245] = v;
	result[246] = v;
	result[247] = v;
	result[248] = v;
	result[249] = v;
	result[250] = v;
	result[251] = v;
	result[252] = v;
	result[253] = v;
	result[254] = v;
	result[255] = v;
end
endmodule

// axi_realigning_burst_reader #(T: type bool #()[32][8], AXI_WIDTH: 256, ADDR_ALIGN: 4, COUNT_TO: 4294967296, ATO: 18446744073709551616)
module axi_realigning_burst_reader_T_type_bool_32_8_AXI_WIDTH_256_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic arvalid,
	input wire arready,
	output /*mux_wire*/ logic[63:0] araddr,
	output /*mux_wire*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[255:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[31:0] count,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic value_valid,
	output /*mux_wire*/ logic[31:0] value[7:0],
	output /*mux_wire*/ logic last
);

/*mux_wire*/ logic _parent_aresetn;
wire _parent_arvalid;
wire[63:0] _parent_araddr;
wire[7:0] _parent_arlen;
wire[2:0] _parent_arsize;
wire[1:0] _parent_arburst;
wire[2:0] _parent_arprot;
wire[3:0] _parent_arcache;
wire[3:0] _parent_arqos;
wire _parent_arlock;
wire[3:0] _parent_arregion;
wire _parent_rready;
/*mux_wire*/ logic _parent_arready;
/*mux_wire*/ logic _parent_rvalid;
/*mux_wire*/ logic[255:0] _parent_rdata;
/*mux_wire*/ logic[1:0] _parent_rresp;
/*mux_wire*/ logic _parent_rlast;
/*mux_wire*/ logic[10:0] _parent_max_in_flight;
wire _parent_may_request_new_burst;
wire[34:0] _22;
assign _22 = count * 4'd8;
/*mux_wire*/ logic _parent_request_new_burst;
/*mux_wire*/ logic[63:0] _parent_start_addr;
/*mux_wire*/ logic[34:0] _parent_count;
/*mux_wire*/ logic _parent_is_ready_to_receive_lots_of_data;
/*state*/ logic[31:0] stored_elements[6:0];
/*state*/ logic[2:0] cur_element_store_align;
wire _parent_element_packet_valid;
wire[31:0] _parent_elements[7:0];
wire[2:0] _parent_chunk_offset;
wire[3:0] _parent_chunk_length;
wire _parent_last;
/*mux_wire*/ logic[31:0] elements[7:0];
/*mux_wire*/ logic[2:0] chunk_offset;
/*mux_wire*/ logic[3:0] chunk_length;
/*mux_wire*/ logic last_2;
/*mux_wire*/ logic[31:0] elements_extended[7:0];
/*mux_wire*/ logic[31:0] rotated_elements[7:0];
wire signed[3:0] _31;
assign _31 = cur_element_store_align - chunk_offset;
wire[2:0] _32;
assign _32 = _31; // == mod 8 (target is 3 bits wide)
/*mux_wire*/ logic[31:0] _RotateRight_data[7:0];
/*mux_wire*/ logic[2:0] _RotateRight_offset;
wire[31:0] _RotateRight_rotated_data[7:0];
/*mux_wire*/ logic[7:0] rotated_strobe;
/*mux_wire*/ logic[2:0] _MakeStrobe_chunk_offset;
/*mux_wire*/ logic[3:0] _MakeStrobe_chunk_length;
wire[7:0] _MakeStrobe_strobe;
/*mux_wire*/ logic[3:0] end_of_element;
wire[3:0] _37;
assign _37 = cur_element_store_align + chunk_length;
wire _39;
assign _39 = end_of_element >= 4'd8;
/*mux_wire*/ logic[255:0] resulting_value_bits;
wire _41;
assign _41 = cur_element_store_align > 1'd0;
wire[31:0] _42 = stored_elements[0];
wire[31:0] _43 = rotated_elements[0];
wire _45;
assign _45 = cur_element_store_align > 1'd1;
wire[31:0] _46 = stored_elements[1];
wire[31:0] _47 = rotated_elements[1];
wire _49;
assign _49 = cur_element_store_align > 2'd2;
wire[31:0] _50 = stored_elements[2];
wire[31:0] _51 = rotated_elements[2];
wire _53;
assign _53 = cur_element_store_align > 2'd3;
wire[31:0] _54 = stored_elements[3];
wire[31:0] _55 = rotated_elements[3];
wire _57;
assign _57 = cur_element_store_align > 3'd4;
wire[31:0] _58 = stored_elements[4];
wire[31:0] _59 = rotated_elements[4];
wire _61;
assign _61 = cur_element_store_align > 3'd5;
wire[31:0] _62 = stored_elements[5];
wire[31:0] _63 = rotated_elements[5];
wire _65;
assign _65 = cur_element_store_align > 3'd6;
wire[31:0] _66 = stored_elements[6];
wire[31:0] _67 = rotated_elements[6];
wire[31:0] _68 = rotated_elements[7];
/*mux_wire*/ logic[255:0] _FromBits_bits;
wire[31:0] _FromBits_value[7:0];
wire[2:0] _73;
assign _73 = end_of_element; // == mod 8 (target is 3 bits wide)
wire _74 = rotated_strobe[0];
wire[31:0] _75 = rotated_elements[0];
wire _76 = rotated_strobe[1];
wire[31:0] _77 = rotated_elements[1];
wire _78 = rotated_strobe[2];
wire[31:0] _79 = rotated_elements[2];
wire _80 = rotated_strobe[3];
wire[31:0] _81 = rotated_elements[3];
wire _82 = rotated_strobe[4];
wire[31:0] _83 = rotated_elements[4];
wire _84 = rotated_strobe[5];
wire[31:0] _85 = rotated_elements[5];
wire _86 = rotated_strobe[6];
wire[31:0] _87 = rotated_elements[6];
wire _89;
assign _89 = !aresetn;
axi_array_burst_reader_AXI_WIDTH_256_ADDR_ALIGN_4_COUNT_TO_34359738368_ATO_18446744073709551616 parent(
	.aclk(aclk),
	.aresetn(_parent_aresetn),
	.arvalid(_parent_arvalid),
	.arready(_parent_arready),
	.araddr(_parent_araddr),
	.arlen(_parent_arlen),
	.arsize(_parent_arsize),
	.arburst(_parent_arburst),
	.arprot(_parent_arprot),
	.arcache(_parent_arcache),
	.arqos(_parent_arqos),
	.arlock(_parent_arlock),
	.arregion(_parent_arregion),
	.rvalid(_parent_rvalid),
	.rready(_parent_rready),
	.rdata(_parent_rdata),
	.rresp(_parent_rresp),
	.rlast(_parent_rlast),
	.is_ready_to_receive_lots_of_data(_parent_is_ready_to_receive_lots_of_data),
	.element_packet_valid(_parent_element_packet_valid),
	.elements(_parent_elements),
	.chunk_offset(_parent_chunk_offset),
	.chunk_length(_parent_chunk_length),
	.last(_parent_last),
	.max_in_flight(_parent_max_in_flight),
	.may_request_new_burst(_parent_may_request_new_burst),
	.request_new_burst(_parent_request_new_burst),
	.start_addr(_parent_start_addr),
	.count(_parent_count)
);
RotateRight_T_type_bool_32_ARRAY_LEN_8 RotateRight(
	.clk(aclk),
	.data(_RotateRight_data),
	.offset(_RotateRight_offset),
	.rotated_data(_RotateRight_rotated_data)
);
MakeStrobe_STROBE_WIDTH_8 MakeStrobe(
	.clk(aclk),
	.chunk_offset(_MakeStrobe_chunk_offset),
	.chunk_length(_MakeStrobe_chunk_length),
	.strobe(_MakeStrobe_strobe)
);
FromBits_T_type_bool_32_8 FromBits(
	.clk(aclk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial _parent_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_aresetn = 1'bx;
	_parent_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_aresetn = _parent_aresetn;
end
always_comb begin // combinatorial arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arvalid = 1'bx;
	arvalid = _parent_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arvalid = arvalid;
end
always_comb begin // combinatorial araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	araddr = 64'dx;
	araddr = _parent_araddr;
end
always_comb begin // combinatorial arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlen = 8'dx;
	arlen = _parent_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = _parent_arsize;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _parent_arburst;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _parent_arprot;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _parent_arcache;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = _parent_arqos;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = _parent_arlock;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = _parent_arregion;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = _parent_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _parent_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_arready = 1'bx;
	_parent_arready = arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_arready = _parent_arready;
end
always_comb begin // combinatorial _parent_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rvalid = 1'bx;
	_parent_rvalid = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rvalid = _parent_rvalid;
end
always_comb begin // combinatorial _parent_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rdata = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_parent_rdata = rdata;
end
always_comb begin // combinatorial _parent_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rresp = 2'bxx;
	_parent_rresp = rresp;
end
always_comb begin // combinatorial _parent_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rlast = 1'bx;
	_parent_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rlast = _parent_rlast;
end
always_comb begin // combinatorial _parent_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_max_in_flight = 11'dx;
	_parent_max_in_flight = max_in_flight;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _parent_may_request_new_burst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial _parent_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_request_new_burst = 1'bx;
	_parent_request_new_burst = 1'b0;
	if(request_new_burst) _parent_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_request_new_burst = _parent_request_new_burst;
end
always_comb begin // combinatorial _parent_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_start_addr = 64'dx;
	if(request_new_burst) _parent_start_addr = start_addr;
end
always_comb begin // combinatorial _parent_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_count = 35'dx;
	if(request_new_burst) _parent_count = _22;
end
always_comb begin // combinatorial _parent_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_is_ready_to_receive_lots_of_data = 1'bx;
	_parent_is_ready_to_receive_lots_of_data = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_is_ready_to_receive_lots_of_data = _parent_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value_valid = 1'bx;
	value_valid = 1'b0;
	if(_parent_element_packet_valid) if(_39) value_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	value_valid = value_valid;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) value[_v0] = _FromBits_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_parent_element_packet_valid) if(_39) last = last_2;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state stored_elements
	if(_parent_element_packet_valid) if(_74) stored_elements[0] <= _75;
	if(_parent_element_packet_valid) if(_76) stored_elements[1] <= _77;
	if(_parent_element_packet_valid) if(_78) stored_elements[2] <= _79;
	if(_parent_element_packet_valid) if(_80) stored_elements[3] <= _81;
	if(_parent_element_packet_valid) if(_82) stored_elements[4] <= _83;
	if(_parent_element_packet_valid) if(_84) stored_elements[5] <= _85;
	if(_parent_element_packet_valid) if(_86) stored_elements[6] <= _87;
end
always_ff @(posedge aclk) begin // state cur_element_store_align
	if(_parent_element_packet_valid) cur_element_store_align <= _73;
	if(_89) cur_element_store_align <= 1'd0;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements[_v0] = _parent_elements[_v0];
end
end
always_comb begin // combinatorial chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_offset = 3'dx;
	if(_parent_element_packet_valid) chunk_offset = _parent_chunk_offset;
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 4'dx;
	if(_parent_element_packet_valid) chunk_length = _parent_chunk_length;
end
always_comb begin // combinatorial last_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last_2 = 1'bx;
	if(_parent_element_packet_valid) last_2 = _parent_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last_2 = last_2;
end
always_comb begin // combinatorial elements_extended
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_extended = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements_extended[_v0] = elements[_v0];
end
end
always_comb begin // combinatorial rotated_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) rotated_elements[_v0] = _RotateRight_rotated_data[_v0];
end
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) _RotateRight_data[_v0] = elements_extended[_v0];
end
end
always_comb begin // combinatorial _RotateRight_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_offset = 3'dx;
	if(_parent_element_packet_valid) _RotateRight_offset = _32;
end
always_comb begin // combinatorial rotated_strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_strobe = 8'bxxxxxxxx;
	if(_parent_element_packet_valid) rotated_strobe = _MakeStrobe_strobe;
end
always_comb begin // combinatorial _MakeStrobe_chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_offset = 3'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_offset = cur_element_store_align;
end
always_comb begin // combinatorial _MakeStrobe_chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_length = 4'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_length = chunk_length;
end
always_comb begin // combinatorial end_of_element
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	end_of_element = 4'dx;
	if(_parent_element_packet_valid) end_of_element = _37;
end
always_comb begin // combinatorial resulting_value_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	resulting_value_bits = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_41) resulting_value_bits[_v0] = _42[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_41) resulting_value_bits[_v0] = _43[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_45) resulting_value_bits[32 + _v0] = _46[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_45) resulting_value_bits[32 + _v0] = _47[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_49) resulting_value_bits[64 + _v0] = _50[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_49) resulting_value_bits[64 + _v0] = _51[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_53) resulting_value_bits[96 + _v0] = _54[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_53) resulting_value_bits[96 + _v0] = _55[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_57) resulting_value_bits[128 + _v0] = _58[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_57) resulting_value_bits[128 + _v0] = _59[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_61) resulting_value_bits[160 + _v0] = _62[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_61) resulting_value_bits[160 + _v0] = _63[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_65) resulting_value_bits[192 + _v0] = _66[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_65) resulting_value_bits[192 + _v0] = _67[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) resulting_value_bits[224 + _v0] = _68[_v0];
end
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_parent_element_packet_valid) if(_39) _FromBits_bits = resulting_value_bits;
end
endmodule

// FromBits #(T: type bool #()[32][8])
module FromBits_T_type_bool_32_8(
	input clk,
	input wire[255:0] bits,
	output /*mux_wire*/ logic[31:0] value[7:0]
);

genvar _g0;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign value[_g0] = bits[(_g0) * 32 +: 32];
end
endgenerate
endmodule

// MakeStrobe #(STROBE_WIDTH: 8)
module MakeStrobe_STROBE_WIDTH_8(
	input clk,
	input wire[2:0] chunk_offset,
	input wire[3:0] chunk_length,
	output /*mux_wire*/ logic[7:0] strobe
);

/*mux_wire*/ logic[7:0] chunk_bits;
wire _2;
assign _2 = chunk_length > 1'd0;
wire _4;
assign _4 = chunk_length > 1'd1;
wire _6;
assign _6 = chunk_length > 2'd2;
wire _8;
assign _8 = chunk_length > 2'd3;
wire _10;
assign _10 = chunk_length > 3'd4;
wire _12;
assign _12 = chunk_length > 3'd5;
wire _14;
assign _14 = chunk_length > 3'd6;
wire _16;
assign _16 = chunk_length > 3'd7;
/*mux_wire*/ logic[7:0] _RotateRight_data;
/*mux_wire*/ logic[2:0] _RotateRight_offset;
wire[7:0] _RotateRight_rotated_data;
RotateRight_T_type_bool_ARRAY_LEN_8 RotateRight(
	.clk(clk),
	.data(_RotateRight_data),
	.offset(_RotateRight_offset),
	.rotated_data(_RotateRight_rotated_data)
);
always_comb begin // combinatorial strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	strobe = 8'bxxxxxxxx;
	strobe = _RotateRight_rotated_data;
end
always_comb begin // combinatorial chunk_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_bits = 8'bxxxxxxxx;
	if(_2) chunk_bits[0] = 1'b1;
	if(!_2) chunk_bits[0] = 1'b0;
	if(_4) chunk_bits[1] = 1'b1;
	if(!_4) chunk_bits[1] = 1'b0;
	if(_6) chunk_bits[2] = 1'b1;
	if(!_6) chunk_bits[2] = 1'b0;
	if(_8) chunk_bits[3] = 1'b1;
	if(!_8) chunk_bits[3] = 1'b0;
	if(_10) chunk_bits[4] = 1'b1;
	if(!_10) chunk_bits[4] = 1'b0;
	if(_12) chunk_bits[5] = 1'b1;
	if(!_12) chunk_bits[5] = 1'b0;
	if(_14) chunk_bits[6] = 1'b1;
	if(!_14) chunk_bits[6] = 1'b0;
	if(_16) chunk_bits[7] = 1'b1;
	if(!_16) chunk_bits[7] = 1'b0;
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = 8'bxxxxxxxx;
	_RotateRight_data = chunk_bits;
end
always_comb begin // combinatorial _RotateRight_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_offset = 3'dx;
	_RotateRight_offset = chunk_offset;
end
endmodule

// RotateRight #(T: type bool #(), ARRAY_LEN: 8)
module RotateRight_T_type_bool_ARRAY_LEN_8(
	input clk,
	input wire[7:0] data,
	input wire[2:0] offset,
	output /*mux_wire*/ logic[7:0] rotated_data
);

/*mux_wire*/ logic[2:0] offset_bits;
/*mux_wire*/ logic[2:0] _UIntToBits_value;
wire[2:0] _UIntToBits_bits;
/*mux_wire*/ logic[7:0] rotate_stages[3:0];
/*mux_wire*/ logic[7:0] from;
wire[7:0] _3 = rotate_stages[0];
wire _4 = offset_bits[0];
wire _5 = from[7];
wire _6 = from[0];
wire _7 = offset_bits[0];
wire _8 = from[0];
wire _9 = from[1];
wire _10 = offset_bits[0];
wire _11 = from[1];
wire _12 = from[2];
wire _13 = offset_bits[0];
wire _14 = from[2];
wire _15 = from[3];
wire _16 = offset_bits[0];
wire _17 = from[3];
wire _18 = from[4];
wire _19 = offset_bits[0];
wire _20 = from[4];
wire _21 = from[5];
wire _22 = offset_bits[0];
wire _23 = from[5];
wire _24 = from[6];
wire _25 = offset_bits[0];
wire _26 = from[6];
wire _27 = from[7];
/*mux_wire*/ logic[7:0] from_2;
wire[7:0] _28 = rotate_stages[1];
wire _29 = offset_bits[1];
wire _30 = from_2[6];
wire _31 = from_2[0];
wire _32 = offset_bits[1];
wire _33 = from_2[7];
wire _34 = from_2[1];
wire _35 = offset_bits[1];
wire _36 = from_2[0];
wire _37 = from_2[2];
wire _38 = offset_bits[1];
wire _39 = from_2[1];
wire _40 = from_2[3];
wire _41 = offset_bits[1];
wire _42 = from_2[2];
wire _43 = from_2[4];
wire _44 = offset_bits[1];
wire _45 = from_2[3];
wire _46 = from_2[5];
wire _47 = offset_bits[1];
wire _48 = from_2[4];
wire _49 = from_2[6];
wire _50 = offset_bits[1];
wire _51 = from_2[5];
wire _52 = from_2[7];
/*mux_wire*/ logic[7:0] from_3;
wire[7:0] _53 = rotate_stages[2];
wire _54 = offset_bits[2];
wire _55 = from_3[4];
wire _56 = from_3[0];
wire _57 = offset_bits[2];
wire _58 = from_3[5];
wire _59 = from_3[1];
wire _60 = offset_bits[2];
wire _61 = from_3[6];
wire _62 = from_3[2];
wire _63 = offset_bits[2];
wire _64 = from_3[7];
wire _65 = from_3[3];
wire _66 = offset_bits[2];
wire _67 = from_3[0];
wire _68 = from_3[4];
wire _69 = offset_bits[2];
wire _70 = from_3[1];
wire _71 = from_3[5];
wire _72 = offset_bits[2];
wire _73 = from_3[2];
wire _74 = from_3[6];
wire _75 = offset_bits[2];
wire _76 = from_3[3];
wire _77 = from_3[7];
wire[7:0] _78 = rotate_stages[3];
UIntToBits_NUM_BITS_3 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = 8'bxxxxxxxx;
	rotated_data = _78;
end
always_comb begin // combinatorial offset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	offset_bits = 3'bxxx;
	offset_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 3'dx;
	_UIntToBits_value = offset;
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{8'bxxxxxxxx, 8'bxxxxxxxx, 8'bxxxxxxxx, 8'bxxxxxxxx};
	rotate_stages[0] = data;
	if(_4) rotate_stages[1][0] = _5;
	if(!_4) rotate_stages[1][0] = _6;
	if(_7) rotate_stages[1][1] = _8;
	if(!_7) rotate_stages[1][1] = _9;
	if(_10) rotate_stages[1][2] = _11;
	if(!_10) rotate_stages[1][2] = _12;
	if(_13) rotate_stages[1][3] = _14;
	if(!_13) rotate_stages[1][3] = _15;
	if(_16) rotate_stages[1][4] = _17;
	if(!_16) rotate_stages[1][4] = _18;
	if(_19) rotate_stages[1][5] = _20;
	if(!_19) rotate_stages[1][5] = _21;
	if(_22) rotate_stages[1][6] = _23;
	if(!_22) rotate_stages[1][6] = _24;
	if(_25) rotate_stages[1][7] = _26;
	if(!_25) rotate_stages[1][7] = _27;
	if(_29) rotate_stages[2][0] = _30;
	if(!_29) rotate_stages[2][0] = _31;
	if(_32) rotate_stages[2][1] = _33;
	if(!_32) rotate_stages[2][1] = _34;
	if(_35) rotate_stages[2][2] = _36;
	if(!_35) rotate_stages[2][2] = _37;
	if(_38) rotate_stages[2][3] = _39;
	if(!_38) rotate_stages[2][3] = _40;
	if(_41) rotate_stages[2][4] = _42;
	if(!_41) rotate_stages[2][4] = _43;
	if(_44) rotate_stages[2][5] = _45;
	if(!_44) rotate_stages[2][5] = _46;
	if(_47) rotate_stages[2][6] = _48;
	if(!_47) rotate_stages[2][6] = _49;
	if(_50) rotate_stages[2][7] = _51;
	if(!_50) rotate_stages[2][7] = _52;
	if(_54) rotate_stages[3][0] = _55;
	if(!_54) rotate_stages[3][0] = _56;
	if(_57) rotate_stages[3][1] = _58;
	if(!_57) rotate_stages[3][1] = _59;
	if(_60) rotate_stages[3][2] = _61;
	if(!_60) rotate_stages[3][2] = _62;
	if(_63) rotate_stages[3][3] = _64;
	if(!_63) rotate_stages[3][3] = _65;
	if(_66) rotate_stages[3][4] = _67;
	if(!_66) rotate_stages[3][4] = _68;
	if(_69) rotate_stages[3][5] = _70;
	if(!_69) rotate_stages[3][5] = _71;
	if(_72) rotate_stages[3][6] = _73;
	if(!_72) rotate_stages[3][6] = _74;
	if(_75) rotate_stages[3][7] = _76;
	if(!_75) rotate_stages[3][7] = _77;
end
always_comb begin // combinatorial from
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from = 8'bxxxxxxxx;
	from = _3;
end
always_comb begin // combinatorial from_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_2 = 8'bxxxxxxxx;
	from_2 = _28;
end
always_comb begin // combinatorial from_3
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_3 = 8'bxxxxxxxx;
	from_3 = _53;
end
endmodule

// RotateRight #(T: type bool #()[32], ARRAY_LEN: 8)
module RotateRight_T_type_bool_32_ARRAY_LEN_8(
	input clk,
	input wire[31:0] data[7:0],
	input wire[2:0] offset,
	output /*mux_wire*/ logic[31:0] rotated_data[7:0]
);

genvar _g0;
/*mux_wire*/ logic[2:0] offset_bits;
/*mux_wire*/ logic[2:0] _UIntToBits_value;
wire[2:0] _UIntToBits_bits;
/*mux_wire*/ logic[31:0] rotate_stages[3:0][7:0];
/*mux_wire*/ logic[31:0] from[7:0];
wire[31:0] _3[7:0];
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _3[_g0] = rotate_stages[0][_g0];
end
endgenerate
wire _4 = offset_bits[0];
wire[31:0] _5 = from[7];
wire[31:0] _6 = from[0];
wire _7 = offset_bits[0];
wire[31:0] _8 = from[0];
wire[31:0] _9 = from[1];
wire _10 = offset_bits[0];
wire[31:0] _11 = from[1];
wire[31:0] _12 = from[2];
wire _13 = offset_bits[0];
wire[31:0] _14 = from[2];
wire[31:0] _15 = from[3];
wire _16 = offset_bits[0];
wire[31:0] _17 = from[3];
wire[31:0] _18 = from[4];
wire _19 = offset_bits[0];
wire[31:0] _20 = from[4];
wire[31:0] _21 = from[5];
wire _22 = offset_bits[0];
wire[31:0] _23 = from[5];
wire[31:0] _24 = from[6];
wire _25 = offset_bits[0];
wire[31:0] _26 = from[6];
wire[31:0] _27 = from[7];
/*mux_wire*/ logic[31:0] from_2[7:0];
wire[31:0] _28[7:0];
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _28[_g0] = rotate_stages[1][_g0];
end
endgenerate
wire _29 = offset_bits[1];
wire[31:0] _30 = from_2[6];
wire[31:0] _31 = from_2[0];
wire _32 = offset_bits[1];
wire[31:0] _33 = from_2[7];
wire[31:0] _34 = from_2[1];
wire _35 = offset_bits[1];
wire[31:0] _36 = from_2[0];
wire[31:0] _37 = from_2[2];
wire _38 = offset_bits[1];
wire[31:0] _39 = from_2[1];
wire[31:0] _40 = from_2[3];
wire _41 = offset_bits[1];
wire[31:0] _42 = from_2[2];
wire[31:0] _43 = from_2[4];
wire _44 = offset_bits[1];
wire[31:0] _45 = from_2[3];
wire[31:0] _46 = from_2[5];
wire _47 = offset_bits[1];
wire[31:0] _48 = from_2[4];
wire[31:0] _49 = from_2[6];
wire _50 = offset_bits[1];
wire[31:0] _51 = from_2[5];
wire[31:0] _52 = from_2[7];
/*mux_wire*/ logic[31:0] from_3[7:0];
wire[31:0] _53[7:0];
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _53[_g0] = rotate_stages[2][_g0];
end
endgenerate
wire _54 = offset_bits[2];
wire[31:0] _55 = from_3[4];
wire[31:0] _56 = from_3[0];
wire _57 = offset_bits[2];
wire[31:0] _58 = from_3[5];
wire[31:0] _59 = from_3[1];
wire _60 = offset_bits[2];
wire[31:0] _61 = from_3[6];
wire[31:0] _62 = from_3[2];
wire _63 = offset_bits[2];
wire[31:0] _64 = from_3[7];
wire[31:0] _65 = from_3[3];
wire _66 = offset_bits[2];
wire[31:0] _67 = from_3[0];
wire[31:0] _68 = from_3[4];
wire _69 = offset_bits[2];
wire[31:0] _70 = from_3[1];
wire[31:0] _71 = from_3[5];
wire _72 = offset_bits[2];
wire[31:0] _73 = from_3[2];
wire[31:0] _74 = from_3[6];
wire _75 = offset_bits[2];
wire[31:0] _76 = from_3[3];
wire[31:0] _77 = from_3[7];
wire[31:0] _78[7:0];
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _78[_g0] = rotate_stages[3][_g0];
end
endgenerate
UIntToBits_NUM_BITS_3 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
rotated_data[_v0] = _78[_v0];
end
end
always_comb begin // combinatorial offset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	offset_bits = 3'bxxx;
	offset_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 3'dx;
	_UIntToBits_value = offset;
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{'{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
rotate_stages[0][_v0] = data[_v0];
end
	if(_4) rotate_stages[1][0] = _5;
	if(!_4) rotate_stages[1][0] = _6;
	if(_7) rotate_stages[1][1] = _8;
	if(!_7) rotate_stages[1][1] = _9;
	if(_10) rotate_stages[1][2] = _11;
	if(!_10) rotate_stages[1][2] = _12;
	if(_13) rotate_stages[1][3] = _14;
	if(!_13) rotate_stages[1][3] = _15;
	if(_16) rotate_stages[1][4] = _17;
	if(!_16) rotate_stages[1][4] = _18;
	if(_19) rotate_stages[1][5] = _20;
	if(!_19) rotate_stages[1][5] = _21;
	if(_22) rotate_stages[1][6] = _23;
	if(!_22) rotate_stages[1][6] = _24;
	if(_25) rotate_stages[1][7] = _26;
	if(!_25) rotate_stages[1][7] = _27;
	if(_29) rotate_stages[2][0] = _30;
	if(!_29) rotate_stages[2][0] = _31;
	if(_32) rotate_stages[2][1] = _33;
	if(!_32) rotate_stages[2][1] = _34;
	if(_35) rotate_stages[2][2] = _36;
	if(!_35) rotate_stages[2][2] = _37;
	if(_38) rotate_stages[2][3] = _39;
	if(!_38) rotate_stages[2][3] = _40;
	if(_41) rotate_stages[2][4] = _42;
	if(!_41) rotate_stages[2][4] = _43;
	if(_44) rotate_stages[2][5] = _45;
	if(!_44) rotate_stages[2][5] = _46;
	if(_47) rotate_stages[2][6] = _48;
	if(!_47) rotate_stages[2][6] = _49;
	if(_50) rotate_stages[2][7] = _51;
	if(!_50) rotate_stages[2][7] = _52;
	if(_54) rotate_stages[3][0] = _55;
	if(!_54) rotate_stages[3][0] = _56;
	if(_57) rotate_stages[3][1] = _58;
	if(!_57) rotate_stages[3][1] = _59;
	if(_60) rotate_stages[3][2] = _61;
	if(!_60) rotate_stages[3][2] = _62;
	if(_63) rotate_stages[3][3] = _64;
	if(!_63) rotate_stages[3][3] = _65;
	if(_66) rotate_stages[3][4] = _67;
	if(!_66) rotate_stages[3][4] = _68;
	if(_69) rotate_stages[3][5] = _70;
	if(!_69) rotate_stages[3][5] = _71;
	if(_72) rotate_stages[3][6] = _73;
	if(!_72) rotate_stages[3][6] = _74;
	if(_75) rotate_stages[3][7] = _76;
	if(!_75) rotate_stages[3][7] = _77;
end
always_comb begin // combinatorial from
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
from[_v0] = _3[_v0];
end
end
always_comb begin // combinatorial from_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_2 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
from_2[_v0] = _28[_v0];
end
end
always_comb begin // combinatorial from_3
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_3 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
from_3[_v0] = _53[_v0];
end
end
endmodule

// axi_array_burst_reader #(AXI_WIDTH: 256, ADDR_ALIGN: 4, COUNT_TO: 34359738368, ATO: 18446744073709551616)
module axi_array_burst_reader_AXI_WIDTH_256_ADDR_ALIGN_4_COUNT_TO_34359738368_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*state*/ logic arvalid,
	input wire arready,
	output /*state*/ logic[63:0] araddr,
	output /*state*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[255:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic element_packet_valid,
	output /*mux_wire*/ logic[31:0] elements[7:0],
	output /*mux_wire*/ logic[2:0] chunk_offset,
	output /*mux_wire*/ logic[3:0] chunk_length,
	output /*mux_wire*/ logic last,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[34:0] count
);

/*latency*/ logic _arvalid_D1; always_ff @(posedge aclk) begin _arvalid_D1 <= arvalid; end
/*latency*/ logic _request_new_burst_D1; always_ff @(posedge aclk) begin _request_new_burst_D1 <= request_new_burst; end
genvar _g0;
localparam[1:0] _1 = 2'b01;
localparam[2:0] _2 = 3'b000;
localparam[3:0] _3 = 4'b0010;
/*mux_wire*/ logic[1:0] _rresp;
/*mux_wire*/ logic _rlast;
/*state*/ logic[11:0] num_in_flight;
/*state*/ logic last_burst_in_flight;
/*mux_wire*/ logic[63:0] next_araddr;
/*latency*/ logic[63:0] _next_araddr_D0; always_ff @(posedge aclk) begin _next_araddr_D0 <= next_araddr; end
wire[58:0] _cur_start_chunk_addr_old;
/*mux_wire*/ logic[58:0] _BitwiseIntConcat_upper;
/*mux_wire*/ logic[4:0] _BitwiseIntConcat_lower;
wire[63:0] _BitwiseIntConcat_v;
/*mux_wire*/ logic[6:0] next_arlen;
/*mux_wire*/ logic next_last_burst_in_flight;
/*latency*/ logic _next_last_burst_in_flight_D0; always_ff @(posedge aclk) begin _next_last_burst_in_flight_D0 <= next_last_burst_in_flight; end
/*mux_wire*/ logic[51:0] cur_burst_addr;
/*mux_wire*/ logic[6:0] cur_align;
/*mux_wire*/ logic[58:0] _BitwiseIntSplit_v;
wire[51:0] _BitwiseIntSplit_upper;
wire[6:0] _BitwiseIntSplit_lower;
/*mux_wire*/ logic chunks_are_left;
/*latency*/ logic _chunks_are_left_D0; always_ff @(posedge aclk) begin _chunks_are_left_D0 <= chunks_are_left; end
wire[32:0] _num_chunks_left_old;
/*latency*/ logic[32:0] __num_chunks_left_old_N1; always_ff @(posedge aclk) begin __num_chunks_left_old_N1 <= _num_chunks_left_old; end
/*latency*/ logic[32:0] __num_chunks_left_old_D0; always_ff @(posedge aclk) begin __num_chunks_left_old_D0 <= __num_chunks_left_old_N1; end
wire _14;
assign _14 = _num_chunks_left_old > 1'd0;
/*latency*/ logic __14_N1; always_ff @(posedge aclk) begin __14_N1 <= _14; end
/*mux_wire*/ logic[6:0] max_chunks_in_this_burst;
/*latency*/ logic[6:0] _max_chunks_in_this_burst_D0; always_ff @(posedge aclk) begin _max_chunks_in_this_burst_D0 <= max_chunks_in_this_burst; end
wire[6:0] _18;
assign _18 = 7'd127 - cur_align;
wire[7:0] _22;
assign _22 = max_chunks_in_this_burst + 1'd1;
wire _23;
assign _23 = __num_chunks_left_old_N1 <= _22;
/*latency*/ logic __23_D0; always_ff @(posedge aclk) begin __23_D0 <= _23; end
/*mux_wire*/ logic[32:0] _IntNarrow_in;
wire[7:0] _IntNarrow_out;
wire[6:0] _26;
assign _26 = _IntNarrow_out - 1'd1;
/*latency*/ logic[6:0] __26_D0; always_ff @(posedge aclk) begin __26_D0 <= _26; end
/*mux_wire*/ logic may_next_arvalid;
/*latency*/ logic _may_next_arvalid_D1; always_ff @(posedge aclk) begin _may_next_arvalid_D1 <= may_next_arvalid; end
wire _num_chunks_left_may_update;
wire _30;
assign _30 = _chunks_are_left_D0 & _num_chunks_left_may_update;
wire _cur_start_chunk_addr_may_update;
wire _32;
assign _32 = _30 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
wire _34;
assign _34 = _32 & _LatencyOffset_out;
wire signed[11:0] _37;
assign _37 = max_in_flight - 8'd128;
wire _38;
assign _38 = $signed({1'b0, num_in_flight}) <= _37;
wire _39;
assign _39 = _34 & _38;
/*mux_wire*/ logic[52:0] next_burst_addr;
wire[52:0] _45;
assign _45 = cur_burst_addr + 1'd1;
/*latency*/ logic[52:0] __45_D0; always_ff @(posedge aclk) begin __45_D0 <= _45; end
/*latency*/ logic[52:0] __45_D1; always_ff @(posedge aclk) begin __45_D1 <= __45_D0; end
/*mux_wire*/ logic[52:0] _BitwiseIntConcat_2_upper;
/*mux_wire*/ logic[6:0] _BitwiseIntConcat_2_lower;
wire[59:0] _BitwiseIntConcat_2_v;
/*mux_wire*/ logic[59:0] _IntNarrow_2_in;
wire[58:0] _IntNarrow_2_out;
/*mux_wire*/ logic _cur_start_chunk_addr_update;
/*mux_wire*/ logic[58:0] _cur_start_chunk_addr_new;
/*mux_wire*/ logic[32:0] next_num_chunks_left;
wire[7:0] _53;
assign _53 = next_arlen + 1'd1;
wire signed[33:0] _54;
assign _54 = __num_chunks_left_old_D0 - _53;
/*mux_wire*/ logic signed[33:0] _IntNarrow_3_in;
wire[32:0] _IntNarrow_3_out;
/*mux_wire*/ logic _num_chunks_left_update;
/*mux_wire*/ logic[32:0] _num_chunks_left_new;
/*mux_wire*/ logic _BoolToInt_i;
wire[0:0] _BoolToInt_o;
wire signed[12:0] _64;
assign _64 = num_in_flight - _BoolToInt_o;
wire _66;
assign _66 = !arvalid;
wire _68;
assign _68 = _66 & may_next_arvalid;
wire[7:0] _71;
assign _71 = next_arlen + 1'd1;
/*mux_wire*/ logic _Ternary_cond;
/*mux_wire*/ logic[7:0] _Ternary_a;
/*mux_wire*/ logic[7:0] _Ternary_b;
wire[7:0] _Ternary_o;
wire signed[12:0] _73;
assign _73 = _64 + $signed({1'b0, _Ternary_o});
/*mux_wire*/ logic signed[12:0] _IntNarrow_4_in;
wire[11:0] _IntNarrow_4_out;
/*state*/ logic[3:0] final_chunk_align;
/*state*/ logic[2:0] cur_chunk_align;
/*mux_wire*/ logic[31:0] elements_2[7:0];
wire[31:0] _75;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _75[_g0] = rdata[_g0];
end
endgenerate
wire[31:0] _76;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _76[_g0] = rdata[32 + _g0];
end
endgenerate
wire[31:0] _77;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _77[_g0] = rdata[64 + _g0];
end
endgenerate
wire[31:0] _78;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _78[_g0] = rdata[96 + _g0];
end
endgenerate
wire[31:0] _79;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _79[_g0] = rdata[128 + _g0];
end
endgenerate
wire[31:0] _80;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _80[_g0] = rdata[160 + _g0];
end
endgenerate
wire[31:0] _81;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _81[_g0] = rdata[192 + _g0];
end
endgenerate
wire[31:0] _82;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _82[_g0] = rdata[224 + _g0];
end
endgenerate
/*mux_wire*/ logic[3:0] num_chunk_elements;
/*mux_wire*/ logic is_last;
wire _85;
assign _85 = num_in_flight == 1'd1;
wire _87;
assign _87 = _85 & last_burst_in_flight;
wire signed[4:0] _91;
assign _91 = final_chunk_align - cur_chunk_align;
/*mux_wire*/ logic signed[4:0] _IntNarrow_5_in;
wire[3:0] _IntNarrow_5_out;
wire[3:0] _93;
assign _93 = 4'd8 - cur_chunk_align;
wire _101;
assign _101 = !chunks_are_left;
/*latency*/ logic __101_D0; always_ff @(posedge aclk) begin __101_D0 <= _101; end
wire _103;
assign _103 = __101_D0 & _num_chunks_left_may_update;
wire _105;
assign _105 = _103 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic[58:0] chunk_addr;
/*latency*/ logic[58:0] _chunk_addr_D1; always_ff @(posedge aclk) begin _chunk_addr_D1 <= chunk_addr; end
/*mux_wire*/ logic[2:0] element_in_chunk_align;
wire[61:0] _107;
assign _107 = start_addr / 3'd4;
/*mux_wire*/ logic[61:0] _BitwiseIntSplit_2_v;
wire[58:0] _BitwiseIntSplit_2_upper;
wire[2:0] _BitwiseIntSplit_2_lower;
/*mux_wire*/ logic[32:0] chunk_count_bits;
/*mux_wire*/ logic[2:0] final_alignment;
wire[35:0] _110;
assign _110 = count + element_in_chunk_align;
/*mux_wire*/ logic[35:0] _BitwiseIntSplit_3_v;
wire[32:0] _BitwiseIntSplit_3_upper;
wire[2:0] _BitwiseIntSplit_3_lower;
/*mux_wire*/ logic[32:0] num_chunks;
/*mux_wire*/ logic is_no_chunks;
wire _113;
assign _113 = chunk_count_bits == 1'd0;
wire _119;
assign _119 = final_alignment != 1'd0;
/*mux_wire*/ logic _BoolToInt_2_i;
wire[0:0] _BoolToInt_2_o;
wire[32:0] _120;
assign _120 = chunk_count_bits + _BoolToInt_2_o;
wire _126;
assign _126 = !is_no_chunks;
wire _129;
assign _129 = final_alignment == 1'd0;
wire _130;
assign _130 = _126 & _129;
/*mux_wire*/ logic _BoolToInt_3_i;
wire[0:0] _BoolToInt_3_o;
/*mux_wire*/ logic[0:0] _BitwiseIntConcat_3_upper;
/*mux_wire*/ logic[2:0] _BitwiseIntConcat_3_lower;
wire[3:0] _BitwiseIntConcat_3_v;
wire _134;
assign _134 = !aresetn;
/*mux_wire*/ logic _cur_start_chunk_addr_rst;
wire _136;
assign _136 = !aresetn;
/*mux_wire*/ logic _num_chunks_left_rst;
wire _138;
assign _138 = !aresetn;
SlowState_T_type_int_FROM_0_TO_576460752303423488_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1 cur_start_chunk_addr(
	.clk(aclk),
	.rst(_cur_start_chunk_addr_rst),
	.old(_cur_start_chunk_addr_old),
	.may_update(_cur_start_chunk_addr_may_update),
	.update(_cur_start_chunk_addr_update),
	.new_1(_cur_start_chunk_addr_new)
);
SlowState_T_type_int_FROM_0_TO_4294967299_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0 num_chunks_left(
	.clk(aclk),
	.rst(_num_chunks_left_rst),
	.old(_num_chunks_left_old),
	.may_update(_num_chunks_left_may_update),
	.update(_num_chunks_left_update),
	.new_1(_num_chunks_left_new)
);
BitwiseIntConcat_UPPER_TO_576460752303423488_LOWER_BITS_5 BitwiseIntConcat(
	.clk(aclk),
	.upper(_BitwiseIntConcat_upper),
	.lower(_BitwiseIntConcat_lower),
	.v(_BitwiseIntConcat_v)
);
BitwiseIntSplit_TO_576460752303423488_LOWER_BITS_7 BitwiseIntSplit(
	.clk(aclk),
	.v(_BitwiseIntSplit_v),
	.upper(_BitwiseIntSplit_upper),
	.lower(_BitwiseIntSplit_lower)
);
IntNarrow_FROM_I_0_TO_I_4294967299_FROM_1_TO_129 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
LatencyOffset_T_type_bool_OFFSET_256 LatencyOffset(
	.clk(aclk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
BitwiseIntConcat_UPPER_TO_4503599627370497_LOWER_BITS_7 BitwiseIntConcat_2(
	.clk(aclk),
	.upper(_BitwiseIntConcat_2_upper),
	.lower(_BitwiseIntConcat_2_lower),
	.v(_BitwiseIntConcat_2_v)
);
IntNarrow_FROM_I_0_TO_I_576460752303423616_FROM_0_TO_576460752303423488 IntNarrow_2(
	.clk(aclk),
	.in(_IntNarrow_2_in),
	.out(_IntNarrow_2_out)
);
IntNarrow_FROM_I_128_TO_I_4294967298_FROM_0_TO_4294967299 IntNarrow_3(
	.clk(aclk),
	.in(_IntNarrow_3_in),
	.out(_IntNarrow_3_out)
);
BoolToInt BoolToInt(
	.clk(aclk),
	.i(_BoolToInt_i),
	.o(_BoolToInt_o)
);
Ternary_T_type_int_FROM_0_TO_129 Ternary(
	.clk(aclk),
	.cond(_Ternary_cond),
	.a(_Ternary_a),
	.b(_Ternary_b),
	.o(_Ternary_o)
);
IntNarrow_FROM_I_1_TO_I_3384_FROM_0_TO_3256 IntNarrow_4(
	.clk(aclk),
	.in(_IntNarrow_4_in),
	.out(_IntNarrow_4_out)
);
IntNarrow_FROM_I_7_TO_I_16_FROM_0_TO_9 IntNarrow_5(
	.clk(aclk),
	.in(_IntNarrow_5_in),
	.out(_IntNarrow_5_out)
);
BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_3 BitwiseIntSplit_2(
	.clk(aclk),
	.v(_BitwiseIntSplit_2_v),
	.upper(_BitwiseIntSplit_2_upper),
	.lower(_BitwiseIntSplit_2_lower)
);
BitwiseIntSplit_TO_34359738375_LOWER_BITS_3 BitwiseIntSplit_3(
	.clk(aclk),
	.v(_BitwiseIntSplit_3_v),
	.upper(_BitwiseIntSplit_3_upper),
	.lower(_BitwiseIntSplit_3_lower)
);
BoolToInt BoolToInt_2(
	.clk(aclk),
	.i(_BoolToInt_2_i),
	.o(_BoolToInt_2_o)
);
BoolToInt BoolToInt_3(
	.clk(aclk),
	.i(_BoolToInt_3_i),
	.o(_BoolToInt_3_o)
);
BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_3 BitwiseIntConcat_3(
	.clk(aclk),
	.upper(_BitwiseIntConcat_3_upper),
	.lower(_BitwiseIntConcat_3_lower),
	.v(_BitwiseIntConcat_3_v)
);
always_ff @(posedge aclk) begin // state arvalid
	if(arvalid) if(arready) arvalid <= 1'b0;
	if(!arvalid) if(may_next_arvalid) arvalid <= 1'b1;
	if(_138) arvalid <= 1'b0;
end
always_ff @(posedge aclk) begin // state araddr
	if(!arvalid) if(may_next_arvalid) araddr <= _next_araddr_D0;
end
always_ff @(posedge aclk) begin // state arlen
	if(!arvalid) if(may_next_arvalid) arlen <= next_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = 3'd5;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _1;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _2;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _3;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = 1'd0;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = 1'd0;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rresp = 2'bxx;
	_rresp = rresp;
end
always_comb begin // combinatorial _rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rlast = 1'bx;
	_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_rlast = _rlast;
end
always_comb begin // combinatorial element_packet_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_packet_valid = 1'bx;
	element_packet_valid = 1'b0;
	if(rvalid) element_packet_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	element_packet_valid = element_packet_valid;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(rvalid) elements[_v0] = elements_2[_v0];
end
end
always_comb begin // combinatorial chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_offset = 3'dx;
	if(rvalid) chunk_offset = cur_chunk_align;
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 4'dx;
	if(rvalid) chunk_length = num_chunk_elements;
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(rvalid) last = is_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state num_in_flight
	num_in_flight <= _IntNarrow_4_out;
	if(_138) num_in_flight <= 1'd0;
end
always_ff @(posedge aclk) begin // state last_burst_in_flight
	if(!arvalid) if(may_next_arvalid) last_burst_in_flight <= _next_last_burst_in_flight_D0;
end
always_comb begin // combinatorial next_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_araddr = 64'dx;
	next_araddr = _BitwiseIntConcat_v;
end
always_comb begin // combinatorial _BitwiseIntConcat_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_upper = 59'dx;
	_BitwiseIntConcat_upper = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial _BitwiseIntConcat_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_lower = 5'dx;
	_BitwiseIntConcat_lower = 1'd0;
end
always_comb begin // combinatorial next_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_arlen = 7'dx;
	if(_chunks_are_left_D0) if(__23_D0) next_arlen = __26_D0;
	if(_chunks_are_left_D0) if(!__23_D0) next_arlen = _max_chunks_in_this_burst_D0;
end
always_comb begin // combinatorial next_last_burst_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_last_burst_in_flight = 1'bx;
	next_last_burst_in_flight = 1'b0;
	if(chunks_are_left) if(_23) next_last_burst_in_flight = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	next_last_burst_in_flight = next_last_burst_in_flight;
end
always_comb begin // combinatorial cur_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_burst_addr = 52'dx;
	cur_burst_addr = _BitwiseIntSplit_upper;
end
always_comb begin // combinatorial cur_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_align = 7'dx;
	cur_align = _BitwiseIntSplit_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_v = 59'dx;
	_BitwiseIntSplit_v = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial chunks_are_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunks_are_left = 1'bx;
	chunks_are_left = __14_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunks_are_left = chunks_are_left;
end
always_comb begin // combinatorial max_chunks_in_this_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	max_chunks_in_this_burst = 7'dx;
	if(chunks_are_left) max_chunks_in_this_burst = _18;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 33'dx;
	if(chunks_are_left) if(_23) _IntNarrow_in = __num_chunks_left_old_N1;
end
always_comb begin // combinatorial may_next_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_next_arvalid = 1'bx;
	may_next_arvalid = _39;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_next_arvalid = may_next_arvalid;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial next_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_burst_addr = 53'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) next_burst_addr = __45_D1;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_upper = 53'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_upper = next_burst_addr;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_lower = 7'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_lower = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_2_in = 60'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _IntNarrow_2_in = _BitwiseIntConcat_2_v;
end
always_comb begin // combinatorial _cur_start_chunk_addr_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_update = 1'bx;
	_cur_start_chunk_addr_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _cur_start_chunk_addr_update = 1'b1;
	if(request_new_burst) _cur_start_chunk_addr_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_update = _cur_start_chunk_addr_update;
end
always_comb begin // combinatorial _cur_start_chunk_addr_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_new = 59'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _cur_start_chunk_addr_new = _IntNarrow_2_out;
	if(_request_new_burst_D1) _cur_start_chunk_addr_new = _chunk_addr_D1;
end
always_comb begin // combinatorial next_num_chunks_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_num_chunks_left = 33'dx;
	if(!arvalid) if(may_next_arvalid) next_num_chunks_left = _IntNarrow_3_out;
end
always_comb begin // combinatorial _IntNarrow_3_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_3_in = 34'sdx;
	if(!arvalid) if(may_next_arvalid) _IntNarrow_3_in = _54;
end
always_comb begin // combinatorial _num_chunks_left_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_update = 1'bx;
	_num_chunks_left_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_update = 1'b1;
	if(request_new_burst) _num_chunks_left_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_update = _num_chunks_left_update;
end
always_comb begin // combinatorial _num_chunks_left_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_new = 33'dx;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_new = next_num_chunks_left;
	if(request_new_burst) _num_chunks_left_new = num_chunks;
end
always_comb begin // combinatorial _BoolToInt_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_i = 1'bx;
	_BoolToInt_i = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_i = _BoolToInt_i;
end
always_comb begin // combinatorial _Ternary_cond
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_cond = 1'bx;
	_Ternary_cond = _68;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Ternary_cond = _Ternary_cond;
end
always_comb begin // combinatorial _Ternary_a
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_a = 8'dx;
	_Ternary_a = _71;
end
always_comb begin // combinatorial _Ternary_b
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_b = 8'dx;
	_Ternary_b = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_4_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_4_in = 13'sdx;
	_IntNarrow_4_in = _73;
end
always_ff @(posedge aclk) begin // state final_chunk_align
	if(request_new_burst) final_chunk_align <= _BitwiseIntConcat_3_v;
end
always_ff @(posedge aclk) begin // state cur_chunk_align
	if(rvalid) cur_chunk_align <= 1'd0;
	if(request_new_burst) cur_chunk_align <= element_in_chunk_align;
end
always_comb begin // combinatorial elements_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_2 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	if(rvalid) elements_2[0] = _75;
	if(rvalid) elements_2[1] = _76;
	if(rvalid) elements_2[2] = _77;
	if(rvalid) elements_2[3] = _78;
	if(rvalid) elements_2[4] = _79;
	if(rvalid) elements_2[5] = _80;
	if(rvalid) elements_2[6] = _81;
	if(rvalid) elements_2[7] = _82;
end
always_comb begin // combinatorial num_chunk_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunk_elements = 4'dx;
	if(rvalid) if(is_last) num_chunk_elements = _IntNarrow_5_out;
	if(rvalid) if(!is_last) num_chunk_elements = _93;
end
always_comb begin // combinatorial is_last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_last = 1'bx;
	if(rvalid) is_last = _87;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_last = is_last;
end
always_comb begin // combinatorial _IntNarrow_5_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_5_in = 5'sdx;
	if(rvalid) if(is_last) _IntNarrow_5_in = _91;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _105;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial chunk_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_addr = 59'dx;
	if(request_new_burst) chunk_addr = _BitwiseIntSplit_2_upper;
end
always_comb begin // combinatorial element_in_chunk_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_in_chunk_align = 3'dx;
	if(request_new_burst) element_in_chunk_align = _BitwiseIntSplit_2_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_2_v = 62'dx;
	if(request_new_burst) _BitwiseIntSplit_2_v = _107;
end
always_comb begin // combinatorial chunk_count_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_count_bits = 33'dx;
	if(request_new_burst) chunk_count_bits = _BitwiseIntSplit_3_upper;
end
always_comb begin // combinatorial final_alignment
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	final_alignment = 3'dx;
	if(request_new_burst) final_alignment = _BitwiseIntSplit_3_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_3_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_3_v = 36'dx;
	if(request_new_burst) _BitwiseIntSplit_3_v = _110;
end
always_comb begin // combinatorial num_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunks = 33'dx;
	if(request_new_burst) if(is_no_chunks) num_chunks = 1'd1;
	if(request_new_burst) if(!is_no_chunks) num_chunks = _120;
end
always_comb begin // combinatorial is_no_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_no_chunks = 1'bx;
	if(request_new_burst) is_no_chunks = _113;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_no_chunks = is_no_chunks;
end
always_comb begin // combinatorial _BoolToInt_2_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_2_i = 1'bx;
	if(request_new_burst) if(!is_no_chunks) _BoolToInt_2_i = _119;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_2_i = _BoolToInt_2_i;
end
always_comb begin // combinatorial _BoolToInt_3_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_3_i = 1'bx;
	if(request_new_burst) _BoolToInt_3_i = _130;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_3_i = _BoolToInt_3_i;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_upper = 1'dx;
	if(request_new_burst) _BitwiseIntConcat_3_upper = _BoolToInt_3_o;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BitwiseIntConcat_3_upper = _BitwiseIntConcat_3_upper;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_lower = 3'dx;
	if(request_new_burst) _BitwiseIntConcat_3_lower = final_alignment;
end
always_comb begin // combinatorial _cur_start_chunk_addr_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_rst = 1'bx;
	_cur_start_chunk_addr_rst = _134;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_rst = _cur_start_chunk_addr_rst;
end
always_comb begin // combinatorial _num_chunks_left_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_rst = 1'bx;
	_num_chunks_left_rst = _136;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_rst = _num_chunks_left_rst;
end
endmodule

// BitwiseIntConcat #(UPPER_TO: 2, LOWER_BITS: 3)
module BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_3(
	input clk,
	input wire[0:0] upper,
	input wire[2:0] lower,
	output /*mux_wire*/ logic[3:0] v
);

/*mux_wire*/ logic[3:0] v_bits;
/*mux_wire*/ logic[2:0] _UIntToBits_value;
wire[2:0] _UIntToBits_bits;
/*mux_wire*/ logic[0:0] _UIntToBits_2_value;
wire[0:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[3:0] _FromBits_bits;
wire[3:0] _FromBits_value;
UIntToBits_NUM_BITS_3 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_1 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_16 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 4'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 4'bxxxx;
	for(int _v0 = 0; _v0 < 3; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
v_bits[3 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 3'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 1'dx;
	_UIntToBits_2_value = upper;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_UIntToBits_2_value = _UIntToBits_2_value;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 4'bxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 16))
module FromBits_T_type_int_FROM_0_TO_16(
	input clk,
	input wire[3:0] bits,
	output /*mux_wire*/ logic[3:0] value
);

assign value = bits;
endmodule

// BitwiseIntSplit #(TO: 34359738375, LOWER_BITS: 3)
module BitwiseIntSplit_TO_34359738375_LOWER_BITS_3(
	input clk,
	input wire[35:0] v,
	output /*mux_wire*/ logic[32:0] upper,
	output /*mux_wire*/ logic[2:0] lower
);

genvar _g0;
/*mux_wire*/ logic[35:0] v_bits;
/*mux_wire*/ logic[35:0] _UIntToBits_value;
wire[35:0] _UIntToBits_bits;
wire[2:0] _2;
generate
for(_g0 = 0; _g0 < 3; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[2:0] _BitsToUInt_bits;
wire[2:0] _BitsToUInt_value;
wire[32:0] _3;
generate
for(_g0 = 0; _g0 < 33; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[3 + _g0];
end
endgenerate
/*mux_wire*/ logic[32:0] _FromBits_bits;
wire[32:0] _FromBits_value;
UIntToBits_NUM_BITS_36 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_3 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_4294967297 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 33'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 3'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 36'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 36'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 3'bxxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// UIntToBits #(NUM_BITS: 36)
module UIntToBits_NUM_BITS_36(
	input clk,
	input wire[35:0] value,
	output /*mux_wire*/ logic[35:0] bits
);

	assign bits = value;
endmodule

// BitwiseIntSplit #(TO: 4611686018427387904, LOWER_BITS: 3)
module BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_3(
	input clk,
	input wire[61:0] v,
	output /*mux_wire*/ logic[58:0] upper,
	output /*mux_wire*/ logic[2:0] lower
);

genvar _g0;
/*mux_wire*/ logic[61:0] v_bits;
/*mux_wire*/ logic[61:0] _UIntToBits_value;
wire[61:0] _UIntToBits_bits;
wire[2:0] _2;
generate
for(_g0 = 0; _g0 < 3; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[2:0] _BitsToUInt_bits;
wire[2:0] _BitsToUInt_value;
wire[58:0] _3;
generate
for(_g0 = 0; _g0 < 59; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[3 + _g0];
end
endgenerate
/*mux_wire*/ logic[58:0] _FromBits_bits;
wire[58:0] _FromBits_value;
UIntToBits_NUM_BITS_62 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_3 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_576460752303423488 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 59'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 3'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 62'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 62'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 3'bxxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 59'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 576460752303423488))
module FromBits_T_type_int_FROM_0_TO_576460752303423488(
	input clk,
	input wire[58:0] bits,
	output /*mux_wire*/ logic[58:0] value
);

assign value = bits;
endmodule

// BitsToUInt #(NUM_BITS: 3)
module BitsToUInt_NUM_BITS_3(
	input clk,
	input wire[2:0] bits,
	output /*mux_wire*/ logic[2:0] value
);

	assign value = bits;
endmodule

// IntNarrow #(FROM_I: -7, TO_I: 16, FROM: 0, TO: 9)
module IntNarrow_FROM_I_7_TO_I_16_FROM_0_TO_9(
	input clk,
	input wire signed[4:0] in,
	output /*mux_wire*/ logic[3:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: -1, TO_I: 3384, FROM: 0, TO: 3256)
module IntNarrow_FROM_I_1_TO_I_3384_FROM_0_TO_3256(
	input clk,
	input wire signed[12:0] in,
	output /*mux_wire*/ logic[11:0] out
);

	assign out = in;
endmodule

// Ternary #(T: type int #(FROM: 0, TO: 129))
module Ternary_T_type_int_FROM_0_TO_129(
	input clk,
	input wire cond,
	input wire[7:0] a,
	input wire[7:0] b,
	output /*mux_wire*/ logic[7:0] o
);

always_comb begin // combinatorial o
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	o = 8'dx;
	if(cond) o = a;
	if(!cond) o = b;
end
endmodule

// IntNarrow #(FROM_I: -128, TO_I: 4294967298, FROM: 0, TO: 4294967299)
module IntNarrow_FROM_I_128_TO_I_4294967298_FROM_0_TO_4294967299(
	input clk,
	input wire signed[33:0] in,
	output /*mux_wire*/ logic[32:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 576460752303423616, FROM: 0, TO: 576460752303423488)
module IntNarrow_FROM_I_0_TO_I_576460752303423616_FROM_0_TO_576460752303423488(
	input clk,
	input wire[59:0] in,
	output /*mux_wire*/ logic[58:0] out
);

	assign out = in;
endmodule

// BitwiseIntConcat #(UPPER_TO: 4503599627370497, LOWER_BITS: 7)
module BitwiseIntConcat_UPPER_TO_4503599627370497_LOWER_BITS_7(
	input clk,
	input wire[52:0] upper,
	input wire[6:0] lower,
	output /*mux_wire*/ logic[59:0] v
);

/*mux_wire*/ logic[59:0] v_bits;
/*mux_wire*/ logic[6:0] _UIntToBits_value;
wire[6:0] _UIntToBits_bits;
/*mux_wire*/ logic[52:0] _UIntToBits_2_value;
wire[52:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[59:0] _FromBits_bits;
wire[59:0] _FromBits_value;
UIntToBits_NUM_BITS_7 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_53 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_576460752303423616 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 60'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 60'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 7; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 53; _v0 = _v0 + 1) begin
v_bits[7 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 7'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 53'dx;
	_UIntToBits_2_value = upper;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 60'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 576460752303423616))
module FromBits_T_type_int_FROM_0_TO_576460752303423616(
	input clk,
	input wire[59:0] bits,
	output /*mux_wire*/ logic[59:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 7)
module UIntToBits_NUM_BITS_7(
	input clk,
	input wire[6:0] value,
	output /*mux_wire*/ logic[6:0] bits
);

	assign bits = value;
endmodule

// LatencyOffset #(T: type bool #(), OFFSET: 256)
module LatencyOffset_T_type_bool_OFFSET_256(
	input clk,
	input wire in,
	output /*mux_wire*/ logic out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 4294967299, FROM: 1, TO: 129)
module IntNarrow_FROM_I_0_TO_I_4294967299_FROM_1_TO_129(
	input clk,
	input wire[32:0] in,
	output /*mux_wire*/ logic[7:0] out
);

	assign out = in;
endmodule

// BitwiseIntSplit #(TO: 576460752303423488, LOWER_BITS: 7)
module BitwiseIntSplit_TO_576460752303423488_LOWER_BITS_7(
	input clk,
	input wire[58:0] v,
	output /*mux_wire*/ logic[51:0] upper,
	output /*mux_wire*/ logic[6:0] lower
);

genvar _g0;
/*mux_wire*/ logic[58:0] v_bits;
/*mux_wire*/ logic[58:0] _UIntToBits_value;
wire[58:0] _UIntToBits_bits;
wire[6:0] _2;
generate
for(_g0 = 0; _g0 < 7; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[6:0] _BitsToUInt_bits;
wire[6:0] _BitsToUInt_value;
wire[51:0] _3;
generate
for(_g0 = 0; _g0 < 52; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[7 + _g0];
end
endgenerate
/*mux_wire*/ logic[51:0] _FromBits_bits;
wire[51:0] _FromBits_value;
UIntToBits_NUM_BITS_59 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_7 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_4503599627370496 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 52'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 7'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 59'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 59'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 7'bxxxxxxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 52'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// BitsToUInt #(NUM_BITS: 7)
module BitsToUInt_NUM_BITS_7(
	input clk,
	input wire[6:0] bits,
	output /*mux_wire*/ logic[6:0] value
);

	assign value = bits;
endmodule

// BitwiseIntConcat #(UPPER_TO: 576460752303423488, LOWER_BITS: 5)
module BitwiseIntConcat_UPPER_TO_576460752303423488_LOWER_BITS_5(
	input clk,
	input wire[58:0] upper,
	input wire[4:0] lower,
	output /*mux_wire*/ logic[63:0] v
);

/*mux_wire*/ logic[63:0] v_bits;
/*mux_wire*/ logic[4:0] _UIntToBits_value;
wire[4:0] _UIntToBits_bits;
/*mux_wire*/ logic[58:0] _UIntToBits_2_value;
wire[58:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[63:0] _FromBits_bits;
wire[63:0] _FromBits_value;
UIntToBits_NUM_BITS_5 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_59 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_18446744073709551616 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 64'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 5; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 59; _v0 = _v0 + 1) begin
v_bits[5 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 5'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 59'dx;
	_UIntToBits_2_value = upper;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// UIntToBits #(NUM_BITS: 59)
module UIntToBits_NUM_BITS_59(
	input clk,
	input wire[58:0] value,
	output /*mux_wire*/ logic[58:0] bits
);

	assign bits = value;
endmodule

// SlowState #(T: type int #(FROM: 0, TO: 576460752303423488), RESET_TO: 0, OLD_DELAY: 1, NEW_DELAY: 1)
module SlowState_T_type_int_FROM_0_TO_576460752303423488_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1(
	input clk,
	input wire rst,
	output /*state*/ logic[58:0] old,
	output /*mux_wire*/ logic may_update,
	input wire update,
	input wire[58:0] new_1
);

/*latency*/ logic _update_D1; always_ff @(posedge clk) begin _update_D1 <= update; end
genvar _g0;
/*mux_wire*/ logic _cross_rst_in;
/*mux_wire*/ logic[58:0] new_s;
/*mux_wire*/ logic update_s;
/*mux_wire*/ logic update_old;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
/*latency*/ logic __LatencyOffset_out_N1; always_ff @(posedge clk) begin __LatencyOffset_out_N1 <= _LatencyOffset_out; end
/*mux_wire*/ logic[58:0] new_old;
/*mux_wire*/ logic[58:0] _LatencyOffset_2_in;
wire[58:0] _LatencyOffset_2_out;
wire _cross_rst_out;
/*latency*/ logic __cross_rst_out_D0; always_ff @(posedge clk) begin __cross_rst_out_D0 <= _cross_rst_out; end
/*state*/ logic[1:0] cooldown;
wire _8 = cooldown[0];
wire _11;
assign _11 = update_s | __cross_rst_out_D0;
/*mux_wire*/ logic _Repeat_v;
wire[1:0] _Repeat_result;
wire[0:0] _12;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _12[_g0] = cooldown[1 + _g0];
end
endgenerate
CrossDomain_T_type_bool cross_rst(
	.in_clk(clk),
	.in(_cross_rst_in),
	.out(_cross_rst_out)
);
LatencyOffset_T_type_bool_OFFSET_2 LatencyOffset(
	.clk(clk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
LatencyOffset_T_type_int_FROM_0_TO_576460752303423488_OFFSET_2 LatencyOffset_2(
	.clk(clk),
	.in(_LatencyOffset_2_in),
	.out(_LatencyOffset_2_out)
);
Repeat_T_type_bool_SIZE_2 Repeat(
	.clk(clk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
always_comb begin // combinatorial _cross_rst_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_rst_in = 1'bx;
	_cross_rst_in = rst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_rst_in = _cross_rst_in;
end
always_ff @(posedge clk) begin // state old
	if(_cross_rst_out) old <= 59'd0;
	if(!_cross_rst_out) if(update_old) old <= new_old;
end
always_comb begin // combinatorial new_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_s = 59'dx;
	if(_update_D1) new_s = new_1;
end
always_comb begin // combinatorial update_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_s = 1'bx;
	if(update) update_s = 1'b1;
	if(!update) update_s = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_s = update_s;
end
always_comb begin // combinatorial update_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_old = 1'bx;
	update_old = __LatencyOffset_out_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_old = update_old;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = update_s;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial new_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_old = 59'dx;
	new_old = _LatencyOffset_2_out;
end
always_comb begin // combinatorial _LatencyOffset_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_2_in = 59'dx;
	_LatencyOffset_2_in = new_s;
end
always_comb begin // combinatorial may_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_update = 1'bx;
	may_update = _8;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_update = may_update;
end
always_ff @(posedge clk) begin // state cooldown
	if(_11) cooldown <= _Repeat_result;
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(!_11) cooldown[_v0] <= _12[_v0];
end
	if(!_11) cooldown[1] <= 1'b1;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	if(_11) _Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
endmodule

// LatencyOffset #(T: type int #(FROM: 0, TO: 576460752303423488), OFFSET: -2)
module LatencyOffset_T_type_int_FROM_0_TO_576460752303423488_OFFSET_2(
	input clk,
	input wire[58:0] in,
	output /*mux_wire*/ logic[58:0] out
);

	assign out = in;
endmodule

// benchmark_burst_read #(AXI_WIDTH: 128)
module benchmark_burst_read_AXI_WIDTH_128(
	input aclk,
	input wire aresetn,
	input wire[11:0] s_axi_control_awaddr,
	input wire s_axi_control_awvalid,
	output /*mux_wire*/ logic s_axi_control_awready,
	input wire[31:0] s_axi_control_wdata,
	input wire[3:0] s_axi_control_wstrb,
	input wire s_axi_control_wvalid,
	output /*mux_wire*/ logic s_axi_control_wready,
	output /*mux_wire*/ logic[1:0] s_axi_control_bresp,
	output /*mux_wire*/ logic s_axi_control_bvalid,
	input wire s_axi_control_bready,
	input wire[11:0] s_axi_control_araddr,
	input wire s_axi_control_arvalid,
	output /*mux_wire*/ logic s_axi_control_arready,
	output /*mux_wire*/ logic[31:0] s_axi_control_rdata,
	output /*mux_wire*/ logic[1:0] s_axi_control_rresp,
	output /*mux_wire*/ logic s_axi_control_rvalid,
	input wire s_axi_control_rready,
	output /*mux_wire*/ logic m_axi_awvalid,
	input wire m_axi_awready,
	output /*mux_wire*/ logic[63:0] m_axi_awaddr,
	output /*mux_wire*/ logic[7:0] m_axi_awlen,
	output /*mux_wire*/ logic[1:0] m_axi_awburst,
	output /*mux_wire*/ logic[3:0] m_axi_awcache,
	output /*mux_wire*/ logic m_axi_wvalid,
	input wire m_axi_wready,
	output /*mux_wire*/ logic[127:0] m_axi_wdata,
	output /*mux_wire*/ logic[15:0] m_axi_wstrb,
	output /*mux_wire*/ logic m_axi_wlast,
	input wire m_axi_bvalid,
	output /*mux_wire*/ logic m_axi_bready,
	input wire[1:0] m_axi_bresp,
	output /*mux_wire*/ logic m_axi_arvalid,
	input wire m_axi_arready,
	output /*mux_wire*/ logic[63:0] m_axi_araddr,
	output /*mux_wire*/ logic[7:0] m_axi_arlen,
	output /*mux_wire*/ logic[2:0] m_axi_arsize,
	output /*mux_wire*/ logic[1:0] m_axi_arburst,
	input wire m_axi_rvalid,
	output /*mux_wire*/ logic m_axi_rready,
	input wire[127:0] m_axi_rdata,
	input wire[1:0] m_axi_rresp,
	input wire m_axi_rlast,
	output /*mux_wire*/ logic[2:0] m_axi_arprot,
	output /*mux_wire*/ logic[3:0] m_axi_arcache,
	output /*mux_wire*/ logic[3:0] m_axi_arqos,
	output /*mux_wire*/ logic m_axi_arlock,
	output /*mux_wire*/ logic[3:0] m_axi_arregion
);

genvar _g0;
/*mux_wire*/ logic _ctrl_aresetn;
wire _ctrl_awready;
wire _ctrl_wready;
wire[1:0] _ctrl_bresp;
wire _ctrl_bvalid;
wire _ctrl_arready;
wire[31:0] _ctrl_rdata;
wire[1:0] _ctrl_rresp;
wire _ctrl_rvalid;
/*mux_wire*/ logic[11:0] _ctrl_awaddr;
/*mux_wire*/ logic _ctrl_awvalid;
/*mux_wire*/ logic[31:0] _ctrl_wdata;
/*mux_wire*/ logic[3:0] _ctrl_wstrb;
/*mux_wire*/ logic _ctrl_wvalid;
/*mux_wire*/ logic _ctrl_bready;
/*mux_wire*/ logic[11:0] _ctrl_araddr;
/*mux_wire*/ logic _ctrl_arvalid;
/*mux_wire*/ logic _ctrl_rready;
/*mux_wire*/ logic _reader_aresetn;
/*mux_wire*/ logic _writer_aresetn;
wire _writer_awvalid;
wire[63:0] _writer_awaddr;
wire[7:0] _writer_awlen;
wire[1:0] _writer_awburst;
wire[3:0] _writer_awcache;
wire _writer_wvalid;
wire[127:0] _writer_wdata;
wire[15:0] _writer_wstrb;
wire _writer_wlast;
wire _writer_bready;
/*mux_wire*/ logic _writer_awready;
/*mux_wire*/ logic _writer_wready;
/*mux_wire*/ logic _writer_bvalid;
/*mux_wire*/ logic[1:0] _writer_bresp;
wire _reader_arvalid;
wire[63:0] _reader_araddr;
wire[7:0] _reader_arlen;
wire[2:0] _reader_arsize;
wire[1:0] _reader_arburst;
wire _reader_rready;
/*mux_wire*/ logic _reader_arready;
/*mux_wire*/ logic _reader_rvalid;
/*mux_wire*/ logic[127:0] _reader_rdata;
/*mux_wire*/ logic[1:0] _reader_rresp;
/*mux_wire*/ logic _reader_rlast;
/*mux_wire*/ logic[63:0] addr_a_bits;
wire[31:0] _ctrl_input_regs[3:0];
wire[31:0] _46 = _ctrl_input_regs[0];
wire[31:0] _47 = _ctrl_input_regs[1];
/*mux_wire*/ logic[63:0] start_addr;
/*mux_wire*/ logic[63:0] _BitsToUInt_bits;
wire[63:0] _BitsToUInt_value;
/*mux_wire*/ logic[31:0] num_to_transfer;
wire[31:0] _49 = _ctrl_input_regs[2];
/*mux_wire*/ logic[31:0] _BitsToUInt_2_bits;
wire[31:0] _BitsToUInt_2_value;
/*mux_wire*/ logic[31:0] _IntNarrow_in;
wire[31:0] _IntNarrow_out;
/*mux_wire*/ logic[31:0] config_bits;
wire[31:0] _50 = _ctrl_input_regs[3];
wire[2:0] _51;
generate
for(_g0 = 0; _g0 < 3; _g0 = _g0 + 1) begin
assign _51[_g0] = config_bits[5 + _g0];
end
endgenerate
wire[3:0] _52;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _52[_g0] = config_bits[8 + _g0];
end
endgenerate
wire[3:0] _53;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _53[_g0] = config_bits[12 + _g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_3_bits;
wire[3:0] _BitsToUInt_3_value;
wire _54 = config_bits[16];
wire[3:0] _55;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _55[_g0] = config_bits[17 + _g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_4_bits;
wire[3:0] _BitsToUInt_4_value;
wire[10:0] _56;
generate
for(_g0 = 0; _g0 < 11; _g0 = _g0 + 1) begin
assign _56[_g0] = config_bits[21 + _g0];
end
endgenerate
/*mux_wire*/ logic[10:0] _BitsToUInt_5_bits;
wire[10:0] _BitsToUInt_5_value;
/*mux_wire*/ logic[10:0] _reader_max_in_flight;
/*state*/ logic[63:0] cycles_since_reset;
wire[64:0] _59;
assign _59 = cycles_since_reset + 1'd1;
wire[63:0] _60;
assign _60 = _59; // == mod 18446744073709551616 (target is 64 bits wide)
/*mux_wire*/ logic[63:0] cycles_since_reset_bits;
/*mux_wire*/ logic[63:0] _UIntToBits_value;
wire[63:0] _UIntToBits_bits;
/*latency*/ logic[63:0] __UIntToBits_bits_D1; always_ff @(posedge aclk) begin __UIntToBits_bits_D1 <= _UIntToBits_bits; end
/*latency*/ logic[63:0] __UIntToBits_bits_D2; always_ff @(posedge aclk) begin __UIntToBits_bits_D2 <= __UIntToBits_bits_D1; end
/*latency*/ logic[63:0] __UIntToBits_bits_D3; always_ff @(posedge aclk) begin __UIntToBits_bits_D3 <= __UIntToBits_bits_D2; end
/*state*/ logic[63:0] cycles_since_reset_at_start;
/*state*/ logic running;
/*state*/ logic[31:0] num_cycles_running;
/*state*/ logic[31:0] hash;
wire _ctrl_start;
/*latency*/ logic __ctrl_start_D1; always_ff @(posedge aclk) begin __ctrl_start_D1 <= _ctrl_start; end
/*latency*/ logic __ctrl_start_D2; always_ff @(posedge aclk) begin __ctrl_start_D2 <= __ctrl_start_D1; end
/*latency*/ logic __ctrl_start_D3; always_ff @(posedge aclk) begin __ctrl_start_D3 <= __ctrl_start_D2; end
/*mux_wire*/ logic _reader_request_new_burst;
/*mux_wire*/ logic[63:0] _reader_start_addr;
/*mux_wire*/ logic[31:0] _reader_count;
localparam[31:0] _67 = 32'b00000000000000000000000000000000;
wire[32:0] _72;
assign _72 = num_cycles_running + 1'd1;
wire[31:0] _73;
assign _73 = _72; // == mod 4294967296 (target is 32 bits wide)
/*mux_wire*/ logic _reader_is_ready_to_receive_lots_of_data;
wire _reader_value_valid;
/*latency*/ logic __reader_value_valid_D1; always_ff @(posedge aclk) begin __reader_value_valid_D1 <= _reader_value_valid; end
/*latency*/ logic __reader_value_valid_D2; always_ff @(posedge aclk) begin __reader_value_valid_D2 <= __reader_value_valid_D1; end
/*latency*/ logic __reader_value_valid_D3; always_ff @(posedge aclk) begin __reader_value_valid_D3 <= __reader_value_valid_D2; end
wire[31:0] _reader_value[3:0];
wire _reader_last;
/*mux_wire*/ logic[31:0] value[3:0];
/*mux_wire*/ logic last;
/*latency*/ logic _last_D1; always_ff @(posedge aclk) begin _last_D1 <= last; end
/*latency*/ logic _last_D2; always_ff @(posedge aclk) begin _last_D2 <= _last_D1; end
/*latency*/ logic _last_D3; always_ff @(posedge aclk) begin _last_D3 <= _last_D2; end
/*mux_wire*/ logic[31:0] new_hash_contrib;
wire[3:0] _74;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _74[_g0] = value[_g0][0];
end
endgenerate
wire _75;
assign _75 = ^_74;
/*latency*/ logic __75_D1; always_ff @(posedge aclk) begin __75_D1 <= _75; end
/*latency*/ logic __75_D2; always_ff @(posedge aclk) begin __75_D2 <= __75_D1; end
wire[3:0] _76;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _76[_g0] = value[_g0][1];
end
endgenerate
wire _77;
assign _77 = ^_76;
/*latency*/ logic __77_D1; always_ff @(posedge aclk) begin __77_D1 <= _77; end
/*latency*/ logic __77_D2; always_ff @(posedge aclk) begin __77_D2 <= __77_D1; end
wire[3:0] _78;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _78[_g0] = value[_g0][2];
end
endgenerate
wire _79;
assign _79 = ^_78;
/*latency*/ logic __79_D1; always_ff @(posedge aclk) begin __79_D1 <= _79; end
/*latency*/ logic __79_D2; always_ff @(posedge aclk) begin __79_D2 <= __79_D1; end
wire[3:0] _80;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _80[_g0] = value[_g0][3];
end
endgenerate
wire _81;
assign _81 = ^_80;
/*latency*/ logic __81_D1; always_ff @(posedge aclk) begin __81_D1 <= _81; end
/*latency*/ logic __81_D2; always_ff @(posedge aclk) begin __81_D2 <= __81_D1; end
wire[3:0] _82;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _82[_g0] = value[_g0][4];
end
endgenerate
wire _83;
assign _83 = ^_82;
/*latency*/ logic __83_D1; always_ff @(posedge aclk) begin __83_D1 <= _83; end
/*latency*/ logic __83_D2; always_ff @(posedge aclk) begin __83_D2 <= __83_D1; end
wire[3:0] _84;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _84[_g0] = value[_g0][5];
end
endgenerate
wire _85;
assign _85 = ^_84;
/*latency*/ logic __85_D1; always_ff @(posedge aclk) begin __85_D1 <= _85; end
/*latency*/ logic __85_D2; always_ff @(posedge aclk) begin __85_D2 <= __85_D1; end
wire[3:0] _86;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _86[_g0] = value[_g0][6];
end
endgenerate
wire _87;
assign _87 = ^_86;
/*latency*/ logic __87_D1; always_ff @(posedge aclk) begin __87_D1 <= _87; end
/*latency*/ logic __87_D2; always_ff @(posedge aclk) begin __87_D2 <= __87_D1; end
wire[3:0] _88;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _88[_g0] = value[_g0][7];
end
endgenerate
wire _89;
assign _89 = ^_88;
/*latency*/ logic __89_D1; always_ff @(posedge aclk) begin __89_D1 <= _89; end
/*latency*/ logic __89_D2; always_ff @(posedge aclk) begin __89_D2 <= __89_D1; end
wire[3:0] _90;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _90[_g0] = value[_g0][8];
end
endgenerate
wire _91;
assign _91 = ^_90;
/*latency*/ logic __91_D1; always_ff @(posedge aclk) begin __91_D1 <= _91; end
/*latency*/ logic __91_D2; always_ff @(posedge aclk) begin __91_D2 <= __91_D1; end
wire[3:0] _92;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _92[_g0] = value[_g0][9];
end
endgenerate
wire _93;
assign _93 = ^_92;
/*latency*/ logic __93_D1; always_ff @(posedge aclk) begin __93_D1 <= _93; end
/*latency*/ logic __93_D2; always_ff @(posedge aclk) begin __93_D2 <= __93_D1; end
wire[3:0] _94;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _94[_g0] = value[_g0][10];
end
endgenerate
wire _95;
assign _95 = ^_94;
/*latency*/ logic __95_D1; always_ff @(posedge aclk) begin __95_D1 <= _95; end
/*latency*/ logic __95_D2; always_ff @(posedge aclk) begin __95_D2 <= __95_D1; end
wire[3:0] _96;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _96[_g0] = value[_g0][11];
end
endgenerate
wire _97;
assign _97 = ^_96;
/*latency*/ logic __97_D1; always_ff @(posedge aclk) begin __97_D1 <= _97; end
/*latency*/ logic __97_D2; always_ff @(posedge aclk) begin __97_D2 <= __97_D1; end
wire[3:0] _98;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _98[_g0] = value[_g0][12];
end
endgenerate
wire _99;
assign _99 = ^_98;
/*latency*/ logic __99_D1; always_ff @(posedge aclk) begin __99_D1 <= _99; end
/*latency*/ logic __99_D2; always_ff @(posedge aclk) begin __99_D2 <= __99_D1; end
wire[3:0] _100;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _100[_g0] = value[_g0][13];
end
endgenerate
wire _101;
assign _101 = ^_100;
/*latency*/ logic __101_D1; always_ff @(posedge aclk) begin __101_D1 <= _101; end
/*latency*/ logic __101_D2; always_ff @(posedge aclk) begin __101_D2 <= __101_D1; end
wire[3:0] _102;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _102[_g0] = value[_g0][14];
end
endgenerate
wire _103;
assign _103 = ^_102;
/*latency*/ logic __103_D1; always_ff @(posedge aclk) begin __103_D1 <= _103; end
/*latency*/ logic __103_D2; always_ff @(posedge aclk) begin __103_D2 <= __103_D1; end
wire[3:0] _104;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _104[_g0] = value[_g0][15];
end
endgenerate
wire _105;
assign _105 = ^_104;
/*latency*/ logic __105_D1; always_ff @(posedge aclk) begin __105_D1 <= _105; end
/*latency*/ logic __105_D2; always_ff @(posedge aclk) begin __105_D2 <= __105_D1; end
wire[3:0] _106;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _106[_g0] = value[_g0][16];
end
endgenerate
wire _107;
assign _107 = ^_106;
/*latency*/ logic __107_D1; always_ff @(posedge aclk) begin __107_D1 <= _107; end
/*latency*/ logic __107_D2; always_ff @(posedge aclk) begin __107_D2 <= __107_D1; end
wire[3:0] _108;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _108[_g0] = value[_g0][17];
end
endgenerate
wire _109;
assign _109 = ^_108;
/*latency*/ logic __109_D1; always_ff @(posedge aclk) begin __109_D1 <= _109; end
/*latency*/ logic __109_D2; always_ff @(posedge aclk) begin __109_D2 <= __109_D1; end
wire[3:0] _110;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _110[_g0] = value[_g0][18];
end
endgenerate
wire _111;
assign _111 = ^_110;
/*latency*/ logic __111_D1; always_ff @(posedge aclk) begin __111_D1 <= _111; end
/*latency*/ logic __111_D2; always_ff @(posedge aclk) begin __111_D2 <= __111_D1; end
wire[3:0] _112;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _112[_g0] = value[_g0][19];
end
endgenerate
wire _113;
assign _113 = ^_112;
/*latency*/ logic __113_D1; always_ff @(posedge aclk) begin __113_D1 <= _113; end
/*latency*/ logic __113_D2; always_ff @(posedge aclk) begin __113_D2 <= __113_D1; end
wire[3:0] _114;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _114[_g0] = value[_g0][20];
end
endgenerate
wire _115;
assign _115 = ^_114;
/*latency*/ logic __115_D1; always_ff @(posedge aclk) begin __115_D1 <= _115; end
/*latency*/ logic __115_D2; always_ff @(posedge aclk) begin __115_D2 <= __115_D1; end
wire[3:0] _116;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _116[_g0] = value[_g0][21];
end
endgenerate
wire _117;
assign _117 = ^_116;
/*latency*/ logic __117_D1; always_ff @(posedge aclk) begin __117_D1 <= _117; end
/*latency*/ logic __117_D2; always_ff @(posedge aclk) begin __117_D2 <= __117_D1; end
wire[3:0] _118;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _118[_g0] = value[_g0][22];
end
endgenerate
wire _119;
assign _119 = ^_118;
/*latency*/ logic __119_D1; always_ff @(posedge aclk) begin __119_D1 <= _119; end
/*latency*/ logic __119_D2; always_ff @(posedge aclk) begin __119_D2 <= __119_D1; end
wire[3:0] _120;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _120[_g0] = value[_g0][23];
end
endgenerate
wire _121;
assign _121 = ^_120;
/*latency*/ logic __121_D1; always_ff @(posedge aclk) begin __121_D1 <= _121; end
/*latency*/ logic __121_D2; always_ff @(posedge aclk) begin __121_D2 <= __121_D1; end
wire[3:0] _122;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _122[_g0] = value[_g0][24];
end
endgenerate
wire _123;
assign _123 = ^_122;
/*latency*/ logic __123_D1; always_ff @(posedge aclk) begin __123_D1 <= _123; end
/*latency*/ logic __123_D2; always_ff @(posedge aclk) begin __123_D2 <= __123_D1; end
wire[3:0] _124;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _124[_g0] = value[_g0][25];
end
endgenerate
wire _125;
assign _125 = ^_124;
/*latency*/ logic __125_D1; always_ff @(posedge aclk) begin __125_D1 <= _125; end
/*latency*/ logic __125_D2; always_ff @(posedge aclk) begin __125_D2 <= __125_D1; end
wire[3:0] _126;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _126[_g0] = value[_g0][26];
end
endgenerate
wire _127;
assign _127 = ^_126;
/*latency*/ logic __127_D1; always_ff @(posedge aclk) begin __127_D1 <= _127; end
/*latency*/ logic __127_D2; always_ff @(posedge aclk) begin __127_D2 <= __127_D1; end
wire[3:0] _128;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _128[_g0] = value[_g0][27];
end
endgenerate
wire _129;
assign _129 = ^_128;
/*latency*/ logic __129_D1; always_ff @(posedge aclk) begin __129_D1 <= _129; end
/*latency*/ logic __129_D2; always_ff @(posedge aclk) begin __129_D2 <= __129_D1; end
wire[3:0] _130;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _130[_g0] = value[_g0][28];
end
endgenerate
wire _131;
assign _131 = ^_130;
/*latency*/ logic __131_D1; always_ff @(posedge aclk) begin __131_D1 <= _131; end
/*latency*/ logic __131_D2; always_ff @(posedge aclk) begin __131_D2 <= __131_D1; end
wire[3:0] _132;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _132[_g0] = value[_g0][29];
end
endgenerate
wire _133;
assign _133 = ^_132;
/*latency*/ logic __133_D1; always_ff @(posedge aclk) begin __133_D1 <= _133; end
/*latency*/ logic __133_D2; always_ff @(posedge aclk) begin __133_D2 <= __133_D1; end
wire[3:0] _134;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _134[_g0] = value[_g0][30];
end
endgenerate
wire _135;
assign _135 = ^_134;
/*latency*/ logic __135_D1; always_ff @(posedge aclk) begin __135_D1 <= _135; end
/*latency*/ logic __135_D2; always_ff @(posedge aclk) begin __135_D2 <= __135_D1; end
wire[3:0] _136;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _136[_g0] = value[_g0][31];
end
endgenerate
wire _137;
assign _137 = ^_136;
/*latency*/ logic __137_D1; always_ff @(posedge aclk) begin __137_D1 <= _137; end
/*latency*/ logic __137_D2; always_ff @(posedge aclk) begin __137_D2 <= __137_D1; end
/*mux_wire*/ logic[31:0] new_hash;
/*latency*/ logic[31:0] _new_hash_D3; always_ff @(posedge aclk) begin _new_hash_D3 <= new_hash; end
wire[31:0] _140;
assign _140 = hash ^ new_hash_contrib;
/*mux_wire*/ logic[31:0] _UIntToBits_2_value;
wire[31:0] _UIntToBits_2_bits;
/*latency*/ logic[31:0] __UIntToBits_2_bits_D1; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D1 <= _UIntToBits_2_bits; end
/*latency*/ logic[31:0] __UIntToBits_2_bits_D2; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D2 <= __UIntToBits_2_bits_D1; end
/*latency*/ logic[31:0] __UIntToBits_2_bits_D3; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D3 <= __UIntToBits_2_bits_D2; end
wire[31:0] _144;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _144[_g0] = cycles_since_reset_at_start[_g0];
end
endgenerate
wire[31:0] _145;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _145[_g0] = cycles_since_reset_at_start[32 + _g0];
end
endgenerate
wire[31:0] _146;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _146[_g0] = cycles_since_reset_bits[_g0];
end
endgenerate
wire[31:0] _147;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _147[_g0] = cycles_since_reset_bits[32 + _g0];
end
endgenerate
wire[31:0] _148[5:0];
assign _148[0] = __UIntToBits_2_bits_D3;
assign _148[1] = _new_hash_D3;
assign _148[2] = _144;
assign _148[3] = _145;
assign _148[4] = _146;
assign _148[5] = _147;
/*mux_wire*/ logic _ctrl_finish;
/*mux_wire*/ logic[31:0] _ctrl_output_regs[5:0];
wire _153;
assign _153 = !aresetn;
/*latency*/ logic __153_D1; always_ff @(posedge aclk) begin __153_D1 <= _153; end
/*latency*/ logic __153_D2; always_ff @(posedge aclk) begin __153_D2 <= __153_D1; end
localparam[31:0] _155 = 32'b00000000000000000000000000000000;
axi_ctrl_slave_NUM_INPUT_REGS_4_NUM_OUTPUT_REGS_6_ADDR_WIDTH_12_AXI_WIDTH_32 ctrl(
	.aclk(aclk),
	.aresetn(_ctrl_aresetn),
	.awaddr(_ctrl_awaddr),
	.awvalid(_ctrl_awvalid),
	.awready(_ctrl_awready),
	.wdata(_ctrl_wdata),
	.wstrb(_ctrl_wstrb),
	.wvalid(_ctrl_wvalid),
	.wready(_ctrl_wready),
	.bresp(_ctrl_bresp),
	.bvalid(_ctrl_bvalid),
	.bready(_ctrl_bready),
	.araddr(_ctrl_araddr),
	.arvalid(_ctrl_arvalid),
	.arready(_ctrl_arready),
	.rdata(_ctrl_rdata),
	.rresp(_ctrl_rresp),
	.rvalid(_ctrl_rvalid),
	.rready(_ctrl_rready),
	.input_regs(_ctrl_input_regs),
	.start(_ctrl_start),
	.finish(_ctrl_finish),
	.output_regs(_ctrl_output_regs)
);
axi_realigning_burst_reader_T_type_bool_32_4_AXI_WIDTH_128_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616 reader(
	.aclk(aclk),
	.aresetn(_reader_aresetn),
	.arvalid(_reader_arvalid),
	.arready(_reader_arready),
	.araddr(_reader_araddr),
	.arlen(_reader_arlen),
	.arsize(_reader_arsize),
	.arburst(_reader_arburst),
	.arprot(),
	.arcache(),
	.arqos(),
	.arlock(),
	.arregion(),
	.rvalid(_reader_rvalid),
	.rready(_reader_rready),
	.rdata(_reader_rdata),
	.rresp(_reader_rresp),
	.rlast(_reader_rlast),
	.max_in_flight(_reader_max_in_flight),
	.may_request_new_burst(),
	.request_new_burst(_reader_request_new_burst),
	.start_addr(_reader_start_addr),
	.count(_reader_count),
	.is_ready_to_receive_lots_of_data(_reader_is_ready_to_receive_lots_of_data),
	.value_valid(_reader_value_valid),
	.value(_reader_value),
	.last(_reader_last)
);
axi_memory_writer_tie_off_AXI_WIDTH_128 writer(
	.aclk(aclk),
	.aresetn(_writer_aresetn),
	.awvalid(_writer_awvalid),
	.awready(_writer_awready),
	.awaddr(_writer_awaddr),
	.awlen(_writer_awlen),
	.awsize(),
	.awburst(_writer_awburst),
	.awprot(),
	.awcache(_writer_awcache),
	.awqos(),
	.awlock(),
	.awregion(),
	.wvalid(_writer_wvalid),
	.wready(_writer_wready),
	.wdata(_writer_wdata),
	.wstrb(_writer_wstrb),
	.wlast(_writer_wlast),
	.bvalid(_writer_bvalid),
	.bresp(_writer_bresp),
	.bready(_writer_bready)
);
BitsToUInt_NUM_BITS_64 BitsToUInt(
	.clk(aclk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
BitsToUInt_NUM_BITS_32 BitsToUInt_2(
	.clk(aclk),
	.bits(_BitsToUInt_2_bits),
	.value(_BitsToUInt_2_value)
);
IntNarrow_FROM_I_0_TO_I_4294967296_FROM_1_TO_4294967296 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
BitsToUInt_NUM_BITS_4 BitsToUInt_3(
	.clk(aclk),
	.bits(_BitsToUInt_3_bits),
	.value(_BitsToUInt_3_value)
);
BitsToUInt_NUM_BITS_4 BitsToUInt_4(
	.clk(aclk),
	.bits(_BitsToUInt_4_bits),
	.value(_BitsToUInt_4_value)
);
BitsToUInt_NUM_BITS_11 BitsToUInt_5(
	.clk(aclk),
	.bits(_BitsToUInt_5_bits),
	.value(_BitsToUInt_5_value)
);
UIntToBits_NUM_BITS_64 UIntToBits(
	.clk(aclk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_32 UIntToBits_2(
	.clk(aclk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
always_comb begin // combinatorial _ctrl_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_aresetn = 1'bx;
	_ctrl_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_aresetn = _ctrl_aresetn;
end
always_comb begin // combinatorial s_axi_control_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_awready = 1'bx;
	s_axi_control_awready = _ctrl_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_awready = s_axi_control_awready;
end
always_comb begin // combinatorial s_axi_control_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_wready = 1'bx;
	s_axi_control_wready = _ctrl_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_wready = s_axi_control_wready;
end
always_comb begin // combinatorial s_axi_control_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bresp = 2'bxx;
	s_axi_control_bresp = _ctrl_bresp;
end
always_comb begin // combinatorial s_axi_control_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bvalid = 1'bx;
	s_axi_control_bvalid = _ctrl_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_bvalid = s_axi_control_bvalid;
end
always_comb begin // combinatorial s_axi_control_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_arready = 1'bx;
	s_axi_control_arready = _ctrl_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_arready = s_axi_control_arready;
end
always_comb begin // combinatorial s_axi_control_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	s_axi_control_rdata = _ctrl_rdata;
end
always_comb begin // combinatorial s_axi_control_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rresp = 2'bxx;
	s_axi_control_rresp = _ctrl_rresp;
end
always_comb begin // combinatorial s_axi_control_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rvalid = 1'bx;
	s_axi_control_rvalid = _ctrl_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_rvalid = s_axi_control_rvalid;
end
always_comb begin // combinatorial _ctrl_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awaddr = 12'dx;
	_ctrl_awaddr = s_axi_control_awaddr;
end
always_comb begin // combinatorial _ctrl_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awvalid = 1'bx;
	_ctrl_awvalid = s_axi_control_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_awvalid = _ctrl_awvalid;
end
always_comb begin // combinatorial _ctrl_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_ctrl_wdata = s_axi_control_wdata;
end
always_comb begin // combinatorial _ctrl_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wstrb = 4'bxxxx;
	_ctrl_wstrb = s_axi_control_wstrb;
end
always_comb begin // combinatorial _ctrl_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wvalid = 1'bx;
	_ctrl_wvalid = s_axi_control_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_wvalid = _ctrl_wvalid;
end
always_comb begin // combinatorial _ctrl_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_bready = 1'bx;
	_ctrl_bready = s_axi_control_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_bready = _ctrl_bready;
end
always_comb begin // combinatorial _ctrl_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_araddr = 12'dx;
	_ctrl_araddr = s_axi_control_araddr;
end
always_comb begin // combinatorial _ctrl_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_arvalid = 1'bx;
	_ctrl_arvalid = s_axi_control_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_arvalid = _ctrl_arvalid;
end
always_comb begin // combinatorial _ctrl_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_rready = 1'bx;
	_ctrl_rready = s_axi_control_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_rready = _ctrl_rready;
end
always_comb begin // combinatorial _reader_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_aresetn = 1'bx;
	_reader_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_aresetn = _reader_aresetn;
end
always_comb begin // combinatorial _writer_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_aresetn = 1'bx;
	_writer_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_aresetn = _writer_aresetn;
end
always_comb begin // combinatorial m_axi_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awvalid = 1'bx;
	m_axi_awvalid = _writer_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_awvalid = m_axi_awvalid;
end
always_comb begin // combinatorial m_axi_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awaddr = 64'dx;
	m_axi_awaddr = _writer_awaddr;
end
always_comb begin // combinatorial m_axi_awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awlen = 8'dx;
	m_axi_awlen = _writer_awlen;
end
always_comb begin // combinatorial m_axi_awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awburst = 2'bxx;
	m_axi_awburst = _writer_awburst;
end
always_comb begin // combinatorial m_axi_awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awcache = 4'bxxxx;
	m_axi_awcache = _writer_awcache;
end
always_comb begin // combinatorial m_axi_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wvalid = 1'bx;
	m_axi_wvalid = _writer_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wvalid = m_axi_wvalid;
end
always_comb begin // combinatorial m_axi_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wdata = 128'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	m_axi_wdata = _writer_wdata;
end
always_comb begin // combinatorial m_axi_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wstrb = 16'bxxxxxxxxxxxxxxxx;
	m_axi_wstrb = _writer_wstrb;
end
always_comb begin // combinatorial m_axi_wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wlast = 1'bx;
	m_axi_wlast = _writer_wlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wlast = m_axi_wlast;
end
always_comb begin // combinatorial m_axi_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_bready = 1'bx;
	m_axi_bready = _writer_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_bready = m_axi_bready;
end
always_comb begin // combinatorial _writer_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_awready = 1'bx;
	_writer_awready = m_axi_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_awready = _writer_awready;
end
always_comb begin // combinatorial _writer_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_wready = 1'bx;
	_writer_wready = m_axi_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_wready = _writer_wready;
end
always_comb begin // combinatorial _writer_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bvalid = 1'bx;
	_writer_bvalid = m_axi_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_bvalid = _writer_bvalid;
end
always_comb begin // combinatorial _writer_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bresp = 2'bxx;
	_writer_bresp = m_axi_bresp;
end
always_comb begin // combinatorial m_axi_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arvalid = 1'bx;
	m_axi_arvalid = _reader_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arvalid = m_axi_arvalid;
end
always_comb begin // combinatorial m_axi_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_araddr = 64'dx;
	m_axi_araddr = _reader_araddr;
end
always_comb begin // combinatorial m_axi_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlen = 8'dx;
	m_axi_arlen = _reader_arlen;
end
always_comb begin // combinatorial m_axi_arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arsize = 3'dx;
	m_axi_arsize = _reader_arsize;
end
always_comb begin // combinatorial m_axi_arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arburst = 2'bxx;
	m_axi_arburst = _reader_arburst;
end
always_comb begin // combinatorial m_axi_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_rready = 1'bx;
	m_axi_rready = _reader_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_rready = m_axi_rready;
end
always_comb begin // combinatorial _reader_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_arready = 1'bx;
	_reader_arready = m_axi_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_arready = _reader_arready;
end
always_comb begin // combinatorial _reader_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rvalid = 1'bx;
	_reader_rvalid = m_axi_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rvalid = _reader_rvalid;
end
always_comb begin // combinatorial _reader_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rdata = 128'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_reader_rdata = m_axi_rdata;
end
always_comb begin // combinatorial _reader_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rresp = 2'bxx;
	_reader_rresp = m_axi_rresp;
end
always_comb begin // combinatorial _reader_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rlast = 1'bx;
	_reader_rlast = m_axi_rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rlast = _reader_rlast;
end
always_comb begin // combinatorial addr_a_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	addr_a_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[_v0] = _46[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[32 + _v0] = _47[_v0];
end
end
always_comb begin // combinatorial start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	start_addr = 64'dx;
	start_addr = _BitsToUInt_value;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_BitsToUInt_bits = addr_a_bits;
end
always_comb begin // combinatorial num_to_transfer
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_to_transfer = 32'dx;
	num_to_transfer = _IntNarrow_out;
end
always_comb begin // combinatorial _BitsToUInt_2_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_2_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_BitsToUInt_2_bits = _49;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 32'dx;
	_IntNarrow_in = _BitsToUInt_2_value;
end
always_comb begin // combinatorial config_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	config_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	config_bits = _50;
end
always_comb begin // combinatorial m_axi_arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arprot = 3'bxxx;
	m_axi_arprot = _51;
end
always_comb begin // combinatorial m_axi_arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arcache = 4'bxxxx;
	m_axi_arcache = _52;
end
always_comb begin // combinatorial m_axi_arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arqos = 4'dx;
	m_axi_arqos = _BitsToUInt_3_value;
end
always_comb begin // combinatorial _BitsToUInt_3_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_3_bits = 4'bxxxx;
	_BitsToUInt_3_bits = _53;
end
always_comb begin // combinatorial m_axi_arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlock = 1'bx;
	m_axi_arlock = _54;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arlock = m_axi_arlock;
end
always_comb begin // combinatorial m_axi_arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arregion = 4'dx;
	m_axi_arregion = _BitsToUInt_4_value;
end
always_comb begin // combinatorial _BitsToUInt_4_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_4_bits = 4'bxxxx;
	_BitsToUInt_4_bits = _55;
end
always_comb begin // combinatorial _BitsToUInt_5_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_5_bits = 11'bxxxxxxxxxxx;
	_BitsToUInt_5_bits = _56;
end
always_comb begin // combinatorial _reader_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_max_in_flight = 11'dx;
	_reader_max_in_flight = _BitsToUInt_5_value;
end
always_ff @(posedge aclk) begin // state cycles_since_reset
	cycles_since_reset <= _60;
	if(_153) cycles_since_reset <= 1'd0;
end
always_comb begin // combinatorial cycles_since_reset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cycles_since_reset_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	cycles_since_reset_bits = __UIntToBits_bits_D3;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 64'dx;
	_UIntToBits_value = cycles_since_reset;
end
always_ff @(posedge aclk) begin // state cycles_since_reset_at_start
	if(__ctrl_start_D3) cycles_since_reset_at_start <= cycles_since_reset_bits;
end
always_ff @(posedge aclk) begin // state running
	if(_ctrl_start) running <= 1'b1;
	if(_reader_value_valid) if(last) running <= 1'b0;
	if(_153) running <= 1'b0;
end
always_ff @(posedge aclk) begin // state num_cycles_running
	if(_ctrl_start) num_cycles_running <= 1'd0;
	if(running) num_cycles_running <= _73;
	if(_153) num_cycles_running <= 1'd0;
end
always_ff @(posedge aclk) begin // state hash
	if(__ctrl_start_D2) hash <= _67;
	if(__reader_value_valid_D2) hash <= new_hash;
	if(__153_D2) hash <= _155;
end
always_comb begin // combinatorial _reader_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_request_new_burst = 1'bx;
	_reader_request_new_burst = 1'b0;
	if(_ctrl_start) _reader_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_request_new_burst = _reader_request_new_burst;
end
always_comb begin // combinatorial _reader_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_start_addr = 64'dx;
	if(_ctrl_start) _reader_start_addr = start_addr;
end
always_comb begin // combinatorial _reader_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_count = 32'dx;
	if(_ctrl_start) _reader_count = num_to_transfer;
end
always_comb begin // combinatorial _reader_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_is_ready_to_receive_lots_of_data = 1'bx;
	_reader_is_ready_to_receive_lots_of_data = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_is_ready_to_receive_lots_of_data = _reader_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
if(_reader_value_valid) value[_v0] = _reader_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_reader_value_valid) last = _reader_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_comb begin // combinatorial new_hash_contrib
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_hash_contrib = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(__reader_value_valid_D2) new_hash_contrib[0] = __75_D2;
	if(__reader_value_valid_D2) new_hash_contrib[1] = __77_D2;
	if(__reader_value_valid_D2) new_hash_contrib[2] = __79_D2;
	if(__reader_value_valid_D2) new_hash_contrib[3] = __81_D2;
	if(__reader_value_valid_D2) new_hash_contrib[4] = __83_D2;
	if(__reader_value_valid_D2) new_hash_contrib[5] = __85_D2;
	if(__reader_value_valid_D2) new_hash_contrib[6] = __87_D2;
	if(__reader_value_valid_D2) new_hash_contrib[7] = __89_D2;
	if(__reader_value_valid_D2) new_hash_contrib[8] = __91_D2;
	if(__reader_value_valid_D2) new_hash_contrib[9] = __93_D2;
	if(__reader_value_valid_D2) new_hash_contrib[10] = __95_D2;
	if(__reader_value_valid_D2) new_hash_contrib[11] = __97_D2;
	if(__reader_value_valid_D2) new_hash_contrib[12] = __99_D2;
	if(__reader_value_valid_D2) new_hash_contrib[13] = __101_D2;
	if(__reader_value_valid_D2) new_hash_contrib[14] = __103_D2;
	if(__reader_value_valid_D2) new_hash_contrib[15] = __105_D2;
	if(__reader_value_valid_D2) new_hash_contrib[16] = __107_D2;
	if(__reader_value_valid_D2) new_hash_contrib[17] = __109_D2;
	if(__reader_value_valid_D2) new_hash_contrib[18] = __111_D2;
	if(__reader_value_valid_D2) new_hash_contrib[19] = __113_D2;
	if(__reader_value_valid_D2) new_hash_contrib[20] = __115_D2;
	if(__reader_value_valid_D2) new_hash_contrib[21] = __117_D2;
	if(__reader_value_valid_D2) new_hash_contrib[22] = __119_D2;
	if(__reader_value_valid_D2) new_hash_contrib[23] = __121_D2;
	if(__reader_value_valid_D2) new_hash_contrib[24] = __123_D2;
	if(__reader_value_valid_D2) new_hash_contrib[25] = __125_D2;
	if(__reader_value_valid_D2) new_hash_contrib[26] = __127_D2;
	if(__reader_value_valid_D2) new_hash_contrib[27] = __129_D2;
	if(__reader_value_valid_D2) new_hash_contrib[28] = __131_D2;
	if(__reader_value_valid_D2) new_hash_contrib[29] = __133_D2;
	if(__reader_value_valid_D2) new_hash_contrib[30] = __135_D2;
	if(__reader_value_valid_D2) new_hash_contrib[31] = __137_D2;
end
always_comb begin // combinatorial new_hash
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_hash = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(__reader_value_valid_D2) new_hash = _140;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 32'dx;
	if(_reader_value_valid) if(last) _UIntToBits_2_value = num_cycles_running;
end
always_comb begin // combinatorial _ctrl_finish
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_finish = 1'bx;
	_ctrl_finish = 1'b0;
	if(__reader_value_valid_D3) if(_last_D3) _ctrl_finish = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_finish = _ctrl_finish;
end
always_comb begin // combinatorial _ctrl_output_regs
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_output_regs = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
if(__reader_value_valid_D3) if(_last_D3) _ctrl_output_regs[_v0] = _148[_v0];
end
end
endmodule

// axi_memory_writer_tie_off #(AXI_WIDTH: 128)
module axi_memory_writer_tie_off_AXI_WIDTH_128(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic awvalid,
	input wire awready,
	output /*mux_wire*/ logic[63:0] awaddr,
	output /*mux_wire*/ logic[7:0] awlen,
	output /*mux_wire*/ logic[2:0] awsize,
	output /*mux_wire*/ logic[1:0] awburst,
	output /*mux_wire*/ logic[2:0] awprot,
	output /*mux_wire*/ logic[3:0] awcache,
	output /*mux_wire*/ logic[3:0] awqos,
	output /*mux_wire*/ logic awlock,
	output /*mux_wire*/ logic[3:0] awregion,
	output /*mux_wire*/ logic wvalid,
	input wire wready,
	output /*mux_wire*/ logic[127:0] wdata,
	output /*mux_wire*/ logic[15:0] wstrb,
	output /*mux_wire*/ logic wlast,
	input wire bvalid,
	input wire[1:0] bresp,
	output /*mux_wire*/ logic bready
);

/*mux_wire*/ logic _aresetn;
localparam[1:0] _4 = 2'b00;
localparam[2:0] _5 = 3'b000;
localparam[3:0] _6 = 4'b0000;
/*mux_wire*/ logic _Repeat_v;
wire[127:0] _Repeat_result;
/*mux_wire*/ logic _Repeat_2_v;
wire[15:0] _Repeat_2_result;
/*mux_wire*/ logic _awready;
/*mux_wire*/ logic _wready;
/*mux_wire*/ logic _bvalid;
/*mux_wire*/ logic[1:0] _bresp;
Repeat_T_type_bool_SIZE_128 Repeat(
	.clk(aclk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
Repeat_T_type_bool_SIZE_16 Repeat_2(
	.clk(aclk),
	.v(_Repeat_2_v),
	.result(_Repeat_2_result)
);
always_comb begin // combinatorial _aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_aresetn = 1'bx;
	_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_aresetn = _aresetn;
end
always_comb begin // combinatorial awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awvalid = 1'bx;
	awvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awvalid = awvalid;
end
always_comb begin // combinatorial awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awaddr = 64'dx;
	awaddr = 1'd0;
end
always_comb begin // combinatorial awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlen = 8'dx;
	awlen = 1'd0;
end
always_comb begin // combinatorial awsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awsize = 3'dx;
	awsize = 3'd4;
end
always_comb begin // combinatorial awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awburst = 2'bxx;
	awburst = _4;
end
always_comb begin // combinatorial awprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awprot = 3'bxxx;
	awprot = _5;
end
always_comb begin // combinatorial awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awcache = 4'bxxxx;
	awcache = _6;
end
always_comb begin // combinatorial awqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awqos = 4'dx;
	awqos = 1'd0;
end
always_comb begin // combinatorial awlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlock = 1'bx;
	awlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awlock = awlock;
end
always_comb begin // combinatorial awregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awregion = 4'dx;
	awregion = 1'd0;
end
always_comb begin // combinatorial wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wvalid = 1'bx;
	wvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wvalid = wvalid;
end
always_comb begin // combinatorial wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wdata = 128'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	wdata = _Repeat_result;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	_Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
always_comb begin // combinatorial wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wstrb = 16'bxxxxxxxxxxxxxxxx;
	wstrb = _Repeat_2_result;
end
always_comb begin // combinatorial _Repeat_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_2_v = 1'bx;
	_Repeat_2_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_2_v = _Repeat_2_v;
end
always_comb begin // combinatorial wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wlast = 1'bx;
	wlast = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wlast = wlast;
end
always_comb begin // combinatorial bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	bready = 1'bx;
	bready = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	bready = bready;
end
always_comb begin // combinatorial _awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_awready = 1'bx;
	_awready = awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_awready = _awready;
end
always_comb begin // combinatorial _wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_wready = 1'bx;
	_wready = wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_wready = _wready;
end
always_comb begin // combinatorial _bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_bvalid = 1'bx;
	_bvalid = bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_bvalid = _bvalid;
end
always_comb begin // combinatorial _bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_bresp = 2'bxx;
	_bresp = bresp;
end
endmodule

// Repeat #(T: type bool #(), SIZE: 16)
module Repeat_T_type_bool_SIZE_16(
	input clk,
	input wire v,
	output /*mux_wire*/ logic[15:0] result
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = 16'bxxxxxxxxxxxxxxxx;
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
	result[4] = v;
	result[5] = v;
	result[6] = v;
	result[7] = v;
	result[8] = v;
	result[9] = v;
	result[10] = v;
	result[11] = v;
	result[12] = v;
	result[13] = v;
	result[14] = v;
	result[15] = v;
end
endmodule

// Repeat #(T: type bool #(), SIZE: 128)
module Repeat_T_type_bool_SIZE_128(
	input clk,
	input wire v,
	output /*mux_wire*/ logic[127:0] result
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = 128'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
	result[4] = v;
	result[5] = v;
	result[6] = v;
	result[7] = v;
	result[8] = v;
	result[9] = v;
	result[10] = v;
	result[11] = v;
	result[12] = v;
	result[13] = v;
	result[14] = v;
	result[15] = v;
	result[16] = v;
	result[17] = v;
	result[18] = v;
	result[19] = v;
	result[20] = v;
	result[21] = v;
	result[22] = v;
	result[23] = v;
	result[24] = v;
	result[25] = v;
	result[26] = v;
	result[27] = v;
	result[28] = v;
	result[29] = v;
	result[30] = v;
	result[31] = v;
	result[32] = v;
	result[33] = v;
	result[34] = v;
	result[35] = v;
	result[36] = v;
	result[37] = v;
	result[38] = v;
	result[39] = v;
	result[40] = v;
	result[41] = v;
	result[42] = v;
	result[43] = v;
	result[44] = v;
	result[45] = v;
	result[46] = v;
	result[47] = v;
	result[48] = v;
	result[49] = v;
	result[50] = v;
	result[51] = v;
	result[52] = v;
	result[53] = v;
	result[54] = v;
	result[55] = v;
	result[56] = v;
	result[57] = v;
	result[58] = v;
	result[59] = v;
	result[60] = v;
	result[61] = v;
	result[62] = v;
	result[63] = v;
	result[64] = v;
	result[65] = v;
	result[66] = v;
	result[67] = v;
	result[68] = v;
	result[69] = v;
	result[70] = v;
	result[71] = v;
	result[72] = v;
	result[73] = v;
	result[74] = v;
	result[75] = v;
	result[76] = v;
	result[77] = v;
	result[78] = v;
	result[79] = v;
	result[80] = v;
	result[81] = v;
	result[82] = v;
	result[83] = v;
	result[84] = v;
	result[85] = v;
	result[86] = v;
	result[87] = v;
	result[88] = v;
	result[89] = v;
	result[90] = v;
	result[91] = v;
	result[92] = v;
	result[93] = v;
	result[94] = v;
	result[95] = v;
	result[96] = v;
	result[97] = v;
	result[98] = v;
	result[99] = v;
	result[100] = v;
	result[101] = v;
	result[102] = v;
	result[103] = v;
	result[104] = v;
	result[105] = v;
	result[106] = v;
	result[107] = v;
	result[108] = v;
	result[109] = v;
	result[110] = v;
	result[111] = v;
	result[112] = v;
	result[113] = v;
	result[114] = v;
	result[115] = v;
	result[116] = v;
	result[117] = v;
	result[118] = v;
	result[119] = v;
	result[120] = v;
	result[121] = v;
	result[122] = v;
	result[123] = v;
	result[124] = v;
	result[125] = v;
	result[126] = v;
	result[127] = v;
end
endmodule

// axi_realigning_burst_reader #(T: type bool #()[32][4], AXI_WIDTH: 128, ADDR_ALIGN: 4, COUNT_TO: 4294967296, ATO: 18446744073709551616)
module axi_realigning_burst_reader_T_type_bool_32_4_AXI_WIDTH_128_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic arvalid,
	input wire arready,
	output /*mux_wire*/ logic[63:0] araddr,
	output /*mux_wire*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[127:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[31:0] count,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic value_valid,
	output /*mux_wire*/ logic[31:0] value[3:0],
	output /*mux_wire*/ logic last
);

/*mux_wire*/ logic _parent_aresetn;
wire _parent_arvalid;
wire[63:0] _parent_araddr;
wire[7:0] _parent_arlen;
wire[2:0] _parent_arsize;
wire[1:0] _parent_arburst;
wire[2:0] _parent_arprot;
wire[3:0] _parent_arcache;
wire[3:0] _parent_arqos;
wire _parent_arlock;
wire[3:0] _parent_arregion;
wire _parent_rready;
/*mux_wire*/ logic _parent_arready;
/*mux_wire*/ logic _parent_rvalid;
/*mux_wire*/ logic[127:0] _parent_rdata;
/*mux_wire*/ logic[1:0] _parent_rresp;
/*mux_wire*/ logic _parent_rlast;
/*mux_wire*/ logic[10:0] _parent_max_in_flight;
wire _parent_may_request_new_burst;
wire[33:0] _22;
assign _22 = count * 3'd4;
/*mux_wire*/ logic _parent_request_new_burst;
/*mux_wire*/ logic[63:0] _parent_start_addr;
/*mux_wire*/ logic[33:0] _parent_count;
/*mux_wire*/ logic _parent_is_ready_to_receive_lots_of_data;
/*state*/ logic[31:0] stored_elements[2:0];
/*state*/ logic[1:0] cur_element_store_align;
wire _parent_element_packet_valid;
wire[31:0] _parent_elements[3:0];
wire[1:0] _parent_chunk_offset;
wire[2:0] _parent_chunk_length;
wire _parent_last;
/*mux_wire*/ logic[31:0] elements[3:0];
/*mux_wire*/ logic[1:0] chunk_offset;
/*mux_wire*/ logic[2:0] chunk_length;
/*mux_wire*/ logic last_2;
/*mux_wire*/ logic[31:0] elements_extended[3:0];
/*mux_wire*/ logic[31:0] rotated_elements[3:0];
wire signed[2:0] _31;
assign _31 = cur_element_store_align - chunk_offset;
wire[1:0] _32;
assign _32 = _31; // == mod 4 (target is 2 bits wide)
/*mux_wire*/ logic[31:0] _RotateRight_data[3:0];
/*mux_wire*/ logic[1:0] _RotateRight_offset;
wire[31:0] _RotateRight_rotated_data[3:0];
/*mux_wire*/ logic[3:0] rotated_strobe;
/*mux_wire*/ logic[1:0] _MakeStrobe_chunk_offset;
/*mux_wire*/ logic[2:0] _MakeStrobe_chunk_length;
wire[3:0] _MakeStrobe_strobe;
/*mux_wire*/ logic[2:0] end_of_element;
wire[2:0] _37;
assign _37 = cur_element_store_align + chunk_length;
wire _39;
assign _39 = end_of_element >= 3'd4;
/*mux_wire*/ logic[127:0] resulting_value_bits;
wire _41;
assign _41 = cur_element_store_align > 1'd0;
wire[31:0] _42 = stored_elements[0];
wire[31:0] _43 = rotated_elements[0];
wire _45;
assign _45 = cur_element_store_align > 1'd1;
wire[31:0] _46 = stored_elements[1];
wire[31:0] _47 = rotated_elements[1];
wire _49;
assign _49 = cur_element_store_align > 2'd2;
wire[31:0] _50 = stored_elements[2];
wire[31:0] _51 = rotated_elements[2];
wire[31:0] _52 = rotated_elements[3];
/*mux_wire*/ logic[127:0] _FromBits_bits;
wire[31:0] _FromBits_value[3:0];
wire[1:0] _57;
assign _57 = end_of_element; // == mod 4 (target is 2 bits wide)
wire _58 = rotated_strobe[0];
wire[31:0] _59 = rotated_elements[0];
wire _60 = rotated_strobe[1];
wire[31:0] _61 = rotated_elements[1];
wire _62 = rotated_strobe[2];
wire[31:0] _63 = rotated_elements[2];
wire _65;
assign _65 = !aresetn;
axi_array_burst_reader_AXI_WIDTH_128_ADDR_ALIGN_4_COUNT_TO_17179869184_ATO_18446744073709551616 parent(
	.aclk(aclk),
	.aresetn(_parent_aresetn),
	.arvalid(_parent_arvalid),
	.arready(_parent_arready),
	.araddr(_parent_araddr),
	.arlen(_parent_arlen),
	.arsize(_parent_arsize),
	.arburst(_parent_arburst),
	.arprot(_parent_arprot),
	.arcache(_parent_arcache),
	.arqos(_parent_arqos),
	.arlock(_parent_arlock),
	.arregion(_parent_arregion),
	.rvalid(_parent_rvalid),
	.rready(_parent_rready),
	.rdata(_parent_rdata),
	.rresp(_parent_rresp),
	.rlast(_parent_rlast),
	.is_ready_to_receive_lots_of_data(_parent_is_ready_to_receive_lots_of_data),
	.element_packet_valid(_parent_element_packet_valid),
	.elements(_parent_elements),
	.chunk_offset(_parent_chunk_offset),
	.chunk_length(_parent_chunk_length),
	.last(_parent_last),
	.max_in_flight(_parent_max_in_flight),
	.may_request_new_burst(_parent_may_request_new_burst),
	.request_new_burst(_parent_request_new_burst),
	.start_addr(_parent_start_addr),
	.count(_parent_count)
);
RotateRight_T_type_bool_32_ARRAY_LEN_4 RotateRight(
	.clk(aclk),
	.data(_RotateRight_data),
	.offset(_RotateRight_offset),
	.rotated_data(_RotateRight_rotated_data)
);
MakeStrobe_STROBE_WIDTH_4 MakeStrobe(
	.clk(aclk),
	.chunk_offset(_MakeStrobe_chunk_offset),
	.chunk_length(_MakeStrobe_chunk_length),
	.strobe(_MakeStrobe_strobe)
);
FromBits_T_type_bool_32_4 FromBits(
	.clk(aclk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial _parent_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_aresetn = 1'bx;
	_parent_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_aresetn = _parent_aresetn;
end
always_comb begin // combinatorial arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arvalid = 1'bx;
	arvalid = _parent_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arvalid = arvalid;
end
always_comb begin // combinatorial araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	araddr = 64'dx;
	araddr = _parent_araddr;
end
always_comb begin // combinatorial arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlen = 8'dx;
	arlen = _parent_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = _parent_arsize;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _parent_arburst;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _parent_arprot;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _parent_arcache;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = _parent_arqos;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = _parent_arlock;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = _parent_arregion;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = _parent_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _parent_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_arready = 1'bx;
	_parent_arready = arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_arready = _parent_arready;
end
always_comb begin // combinatorial _parent_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rvalid = 1'bx;
	_parent_rvalid = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rvalid = _parent_rvalid;
end
always_comb begin // combinatorial _parent_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rdata = 128'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_parent_rdata = rdata;
end
always_comb begin // combinatorial _parent_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rresp = 2'bxx;
	_parent_rresp = rresp;
end
always_comb begin // combinatorial _parent_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rlast = 1'bx;
	_parent_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rlast = _parent_rlast;
end
always_comb begin // combinatorial _parent_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_max_in_flight = 11'dx;
	_parent_max_in_flight = max_in_flight;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _parent_may_request_new_burst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial _parent_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_request_new_burst = 1'bx;
	_parent_request_new_burst = 1'b0;
	if(request_new_burst) _parent_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_request_new_burst = _parent_request_new_burst;
end
always_comb begin // combinatorial _parent_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_start_addr = 64'dx;
	if(request_new_burst) _parent_start_addr = start_addr;
end
always_comb begin // combinatorial _parent_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_count = 34'dx;
	if(request_new_burst) _parent_count = _22;
end
always_comb begin // combinatorial _parent_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_is_ready_to_receive_lots_of_data = 1'bx;
	_parent_is_ready_to_receive_lots_of_data = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_is_ready_to_receive_lots_of_data = _parent_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value_valid = 1'bx;
	value_valid = 1'b0;
	if(_parent_element_packet_valid) if(_39) value_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	value_valid = value_valid;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) value[_v0] = _FromBits_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_parent_element_packet_valid) if(_39) last = last_2;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state stored_elements
	if(_parent_element_packet_valid) if(_58) stored_elements[0] <= _59;
	if(_parent_element_packet_valid) if(_60) stored_elements[1] <= _61;
	if(_parent_element_packet_valid) if(_62) stored_elements[2] <= _63;
end
always_ff @(posedge aclk) begin // state cur_element_store_align
	if(_parent_element_packet_valid) cur_element_store_align <= _57;
	if(_65) cur_element_store_align <= 1'd0;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements[_v0] = _parent_elements[_v0];
end
end
always_comb begin // combinatorial chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_offset = 2'dx;
	if(_parent_element_packet_valid) chunk_offset = _parent_chunk_offset;
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 3'dx;
	if(_parent_element_packet_valid) chunk_length = _parent_chunk_length;
end
always_comb begin // combinatorial last_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last_2 = 1'bx;
	if(_parent_element_packet_valid) last_2 = _parent_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last_2 = last_2;
end
always_comb begin // combinatorial elements_extended
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_extended = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements_extended[_v0] = elements[_v0];
end
end
always_comb begin // combinatorial rotated_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) rotated_elements[_v0] = _RotateRight_rotated_data[_v0];
end
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) _RotateRight_data[_v0] = elements_extended[_v0];
end
end
always_comb begin // combinatorial _RotateRight_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_offset = 2'dx;
	if(_parent_element_packet_valid) _RotateRight_offset = _32;
end
always_comb begin // combinatorial rotated_strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_strobe = 4'bxxxx;
	if(_parent_element_packet_valid) rotated_strobe = _MakeStrobe_strobe;
end
always_comb begin // combinatorial _MakeStrobe_chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_offset = 2'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_offset = cur_element_store_align;
end
always_comb begin // combinatorial _MakeStrobe_chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_length = 3'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_length = chunk_length;
end
always_comb begin // combinatorial end_of_element
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	end_of_element = 3'dx;
	if(_parent_element_packet_valid) end_of_element = _37;
end
always_comb begin // combinatorial resulting_value_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	resulting_value_bits = 128'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_41) resulting_value_bits[_v0] = _42[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_41) resulting_value_bits[_v0] = _43[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_45) resulting_value_bits[32 + _v0] = _46[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_45) resulting_value_bits[32 + _v0] = _47[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_49) resulting_value_bits[64 + _v0] = _50[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_49) resulting_value_bits[64 + _v0] = _51[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) resulting_value_bits[96 + _v0] = _52[_v0];
end
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 128'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_parent_element_packet_valid) if(_39) _FromBits_bits = resulting_value_bits;
end
endmodule

// FromBits #(T: type bool #()[32][4])
module FromBits_T_type_bool_32_4(
	input clk,
	input wire[127:0] bits,
	output /*mux_wire*/ logic[31:0] value[3:0]
);

genvar _g0;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign value[_g0] = bits[(_g0) * 32 +: 32];
end
endgenerate
endmodule

// MakeStrobe #(STROBE_WIDTH: 4)
module MakeStrobe_STROBE_WIDTH_4(
	input clk,
	input wire[1:0] chunk_offset,
	input wire[2:0] chunk_length,
	output /*mux_wire*/ logic[3:0] strobe
);

/*mux_wire*/ logic[3:0] chunk_bits;
wire _2;
assign _2 = chunk_length > 1'd0;
wire _4;
assign _4 = chunk_length > 1'd1;
wire _6;
assign _6 = chunk_length > 2'd2;
wire _8;
assign _8 = chunk_length > 2'd3;
/*mux_wire*/ logic[3:0] _RotateRight_data;
/*mux_wire*/ logic[1:0] _RotateRight_offset;
wire[3:0] _RotateRight_rotated_data;
RotateRight_T_type_bool_ARRAY_LEN_4 RotateRight(
	.clk(clk),
	.data(_RotateRight_data),
	.offset(_RotateRight_offset),
	.rotated_data(_RotateRight_rotated_data)
);
always_comb begin // combinatorial strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	strobe = 4'bxxxx;
	strobe = _RotateRight_rotated_data;
end
always_comb begin // combinatorial chunk_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_bits = 4'bxxxx;
	if(_2) chunk_bits[0] = 1'b1;
	if(!_2) chunk_bits[0] = 1'b0;
	if(_4) chunk_bits[1] = 1'b1;
	if(!_4) chunk_bits[1] = 1'b0;
	if(_6) chunk_bits[2] = 1'b1;
	if(!_6) chunk_bits[2] = 1'b0;
	if(_8) chunk_bits[3] = 1'b1;
	if(!_8) chunk_bits[3] = 1'b0;
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = 4'bxxxx;
	_RotateRight_data = chunk_bits;
end
always_comb begin // combinatorial _RotateRight_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_offset = 2'dx;
	_RotateRight_offset = chunk_offset;
end
endmodule

// RotateRight #(T: type bool #(), ARRAY_LEN: 4)
module RotateRight_T_type_bool_ARRAY_LEN_4(
	input clk,
	input wire[3:0] data,
	input wire[1:0] offset,
	output /*mux_wire*/ logic[3:0] rotated_data
);

/*mux_wire*/ logic[1:0] offset_bits;
/*mux_wire*/ logic[1:0] _UIntToBits_value;
wire[1:0] _UIntToBits_bits;
/*mux_wire*/ logic[3:0] rotate_stages[2:0];
/*mux_wire*/ logic[3:0] from;
wire[3:0] _3 = rotate_stages[0];
wire _4 = offset_bits[0];
wire _5 = from[3];
wire _6 = from[0];
wire _7 = offset_bits[0];
wire _8 = from[0];
wire _9 = from[1];
wire _10 = offset_bits[0];
wire _11 = from[1];
wire _12 = from[2];
wire _13 = offset_bits[0];
wire _14 = from[2];
wire _15 = from[3];
/*mux_wire*/ logic[3:0] from_2;
wire[3:0] _16 = rotate_stages[1];
wire _17 = offset_bits[1];
wire _18 = from_2[2];
wire _19 = from_2[0];
wire _20 = offset_bits[1];
wire _21 = from_2[3];
wire _22 = from_2[1];
wire _23 = offset_bits[1];
wire _24 = from_2[0];
wire _25 = from_2[2];
wire _26 = offset_bits[1];
wire _27 = from_2[1];
wire _28 = from_2[3];
wire[3:0] _29 = rotate_stages[2];
UIntToBits_NUM_BITS_2 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = 4'bxxxx;
	rotated_data = _29;
end
always_comb begin // combinatorial offset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	offset_bits = 2'bxx;
	offset_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 2'dx;
	_UIntToBits_value = offset;
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{4'bxxxx, 4'bxxxx, 4'bxxxx};
	rotate_stages[0] = data;
	if(_4) rotate_stages[1][0] = _5;
	if(!_4) rotate_stages[1][0] = _6;
	if(_7) rotate_stages[1][1] = _8;
	if(!_7) rotate_stages[1][1] = _9;
	if(_10) rotate_stages[1][2] = _11;
	if(!_10) rotate_stages[1][2] = _12;
	if(_13) rotate_stages[1][3] = _14;
	if(!_13) rotate_stages[1][3] = _15;
	if(_17) rotate_stages[2][0] = _18;
	if(!_17) rotate_stages[2][0] = _19;
	if(_20) rotate_stages[2][1] = _21;
	if(!_20) rotate_stages[2][1] = _22;
	if(_23) rotate_stages[2][2] = _24;
	if(!_23) rotate_stages[2][2] = _25;
	if(_26) rotate_stages[2][3] = _27;
	if(!_26) rotate_stages[2][3] = _28;
end
always_comb begin // combinatorial from
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from = 4'bxxxx;
	from = _3;
end
always_comb begin // combinatorial from_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_2 = 4'bxxxx;
	from_2 = _16;
end
endmodule

// RotateRight #(T: type bool #()[32], ARRAY_LEN: 4)
module RotateRight_T_type_bool_32_ARRAY_LEN_4(
	input clk,
	input wire[31:0] data[3:0],
	input wire[1:0] offset,
	output /*mux_wire*/ logic[31:0] rotated_data[3:0]
);

genvar _g0;
/*mux_wire*/ logic[1:0] offset_bits;
/*mux_wire*/ logic[1:0] _UIntToBits_value;
wire[1:0] _UIntToBits_bits;
/*mux_wire*/ logic[31:0] rotate_stages[2:0][3:0];
/*mux_wire*/ logic[31:0] from[3:0];
wire[31:0] _3[3:0];
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _3[_g0] = rotate_stages[0][_g0];
end
endgenerate
wire _4 = offset_bits[0];
wire[31:0] _5 = from[3];
wire[31:0] _6 = from[0];
wire _7 = offset_bits[0];
wire[31:0] _8 = from[0];
wire[31:0] _9 = from[1];
wire _10 = offset_bits[0];
wire[31:0] _11 = from[1];
wire[31:0] _12 = from[2];
wire _13 = offset_bits[0];
wire[31:0] _14 = from[2];
wire[31:0] _15 = from[3];
/*mux_wire*/ logic[31:0] from_2[3:0];
wire[31:0] _16[3:0];
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _16[_g0] = rotate_stages[1][_g0];
end
endgenerate
wire _17 = offset_bits[1];
wire[31:0] _18 = from_2[2];
wire[31:0] _19 = from_2[0];
wire _20 = offset_bits[1];
wire[31:0] _21 = from_2[3];
wire[31:0] _22 = from_2[1];
wire _23 = offset_bits[1];
wire[31:0] _24 = from_2[0];
wire[31:0] _25 = from_2[2];
wire _26 = offset_bits[1];
wire[31:0] _27 = from_2[1];
wire[31:0] _28 = from_2[3];
wire[31:0] _29[3:0];
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _29[_g0] = rotate_stages[2][_g0];
end
endgenerate
UIntToBits_NUM_BITS_2 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
rotated_data[_v0] = _29[_v0];
end
end
always_comb begin // combinatorial offset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	offset_bits = 2'bxx;
	offset_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 2'dx;
	_UIntToBits_value = offset;
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{'{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
rotate_stages[0][_v0] = data[_v0];
end
	if(_4) rotate_stages[1][0] = _5;
	if(!_4) rotate_stages[1][0] = _6;
	if(_7) rotate_stages[1][1] = _8;
	if(!_7) rotate_stages[1][1] = _9;
	if(_10) rotate_stages[1][2] = _11;
	if(!_10) rotate_stages[1][2] = _12;
	if(_13) rotate_stages[1][3] = _14;
	if(!_13) rotate_stages[1][3] = _15;
	if(_17) rotate_stages[2][0] = _18;
	if(!_17) rotate_stages[2][0] = _19;
	if(_20) rotate_stages[2][1] = _21;
	if(!_20) rotate_stages[2][1] = _22;
	if(_23) rotate_stages[2][2] = _24;
	if(!_23) rotate_stages[2][2] = _25;
	if(_26) rotate_stages[2][3] = _27;
	if(!_26) rotate_stages[2][3] = _28;
end
always_comb begin // combinatorial from
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
from[_v0] = _3[_v0];
end
end
always_comb begin // combinatorial from_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_2 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
from_2[_v0] = _16[_v0];
end
end
endmodule

// axi_array_burst_reader #(AXI_WIDTH: 128, ADDR_ALIGN: 4, COUNT_TO: 17179869184, ATO: 18446744073709551616)
module axi_array_burst_reader_AXI_WIDTH_128_ADDR_ALIGN_4_COUNT_TO_17179869184_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*state*/ logic arvalid,
	input wire arready,
	output /*state*/ logic[63:0] araddr,
	output /*state*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[127:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic element_packet_valid,
	output /*mux_wire*/ logic[31:0] elements[3:0],
	output /*mux_wire*/ logic[1:0] chunk_offset,
	output /*mux_wire*/ logic[2:0] chunk_length,
	output /*mux_wire*/ logic last,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[33:0] count
);

/*latency*/ logic _arvalid_D1; always_ff @(posedge aclk) begin _arvalid_D1 <= arvalid; end
/*latency*/ logic _request_new_burst_D1; always_ff @(posedge aclk) begin _request_new_burst_D1 <= request_new_burst; end
genvar _g0;
localparam[1:0] _1 = 2'b01;
localparam[2:0] _2 = 3'b000;
localparam[3:0] _3 = 4'b0010;
/*mux_wire*/ logic[1:0] _rresp;
/*mux_wire*/ logic _rlast;
/*state*/ logic[11:0] num_in_flight;
/*state*/ logic last_burst_in_flight;
/*mux_wire*/ logic[63:0] next_araddr;
/*latency*/ logic[63:0] _next_araddr_D0; always_ff @(posedge aclk) begin _next_araddr_D0 <= next_araddr; end
wire[59:0] _cur_start_chunk_addr_old;
/*mux_wire*/ logic[59:0] _BitwiseIntConcat_upper;
/*mux_wire*/ logic[3:0] _BitwiseIntConcat_lower;
wire[63:0] _BitwiseIntConcat_v;
/*mux_wire*/ logic[7:0] next_arlen;
/*mux_wire*/ logic next_last_burst_in_flight;
/*latency*/ logic _next_last_burst_in_flight_D0; always_ff @(posedge aclk) begin _next_last_burst_in_flight_D0 <= next_last_burst_in_flight; end
/*mux_wire*/ logic[51:0] cur_burst_addr;
/*mux_wire*/ logic[7:0] cur_align;
/*mux_wire*/ logic[59:0] _BitwiseIntSplit_v;
wire[51:0] _BitwiseIntSplit_upper;
wire[7:0] _BitwiseIntSplit_lower;
/*mux_wire*/ logic chunks_are_left;
/*latency*/ logic _chunks_are_left_D0; always_ff @(posedge aclk) begin _chunks_are_left_D0 <= chunks_are_left; end
wire[32:0] _num_chunks_left_old;
/*latency*/ logic[32:0] __num_chunks_left_old_N1; always_ff @(posedge aclk) begin __num_chunks_left_old_N1 <= _num_chunks_left_old; end
/*latency*/ logic[32:0] __num_chunks_left_old_D0; always_ff @(posedge aclk) begin __num_chunks_left_old_D0 <= __num_chunks_left_old_N1; end
wire _14;
assign _14 = _num_chunks_left_old > 1'd0;
/*latency*/ logic __14_N1; always_ff @(posedge aclk) begin __14_N1 <= _14; end
/*mux_wire*/ logic[7:0] max_chunks_in_this_burst;
/*latency*/ logic[7:0] _max_chunks_in_this_burst_D0; always_ff @(posedge aclk) begin _max_chunks_in_this_burst_D0 <= max_chunks_in_this_burst; end
wire[7:0] _18;
assign _18 = 8'd255 - cur_align;
wire[8:0] _22;
assign _22 = max_chunks_in_this_burst + 1'd1;
wire _23;
assign _23 = __num_chunks_left_old_N1 <= _22;
/*latency*/ logic __23_D0; always_ff @(posedge aclk) begin __23_D0 <= _23; end
/*mux_wire*/ logic[32:0] _IntNarrow_in;
wire[8:0] _IntNarrow_out;
wire[7:0] _26;
assign _26 = _IntNarrow_out - 1'd1;
/*latency*/ logic[7:0] __26_D0; always_ff @(posedge aclk) begin __26_D0 <= _26; end
/*mux_wire*/ logic may_next_arvalid;
/*latency*/ logic _may_next_arvalid_D1; always_ff @(posedge aclk) begin _may_next_arvalid_D1 <= may_next_arvalid; end
wire _num_chunks_left_may_update;
wire _30;
assign _30 = _chunks_are_left_D0 & _num_chunks_left_may_update;
wire _cur_start_chunk_addr_may_update;
wire _32;
assign _32 = _30 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
wire _34;
assign _34 = _32 & _LatencyOffset_out;
wire signed[11:0] _37;
assign _37 = max_in_flight - 9'd256;
wire _38;
assign _38 = $signed({1'b0, num_in_flight}) <= _37;
wire _39;
assign _39 = _34 & _38;
/*mux_wire*/ logic[52:0] next_burst_addr;
wire[52:0] _45;
assign _45 = cur_burst_addr + 1'd1;
/*latency*/ logic[52:0] __45_D0; always_ff @(posedge aclk) begin __45_D0 <= _45; end
/*latency*/ logic[52:0] __45_D1; always_ff @(posedge aclk) begin __45_D1 <= __45_D0; end
/*mux_wire*/ logic[52:0] _BitwiseIntConcat_2_upper;
/*mux_wire*/ logic[7:0] _BitwiseIntConcat_2_lower;
wire[60:0] _BitwiseIntConcat_2_v;
/*mux_wire*/ logic[60:0] _IntNarrow_2_in;
wire[59:0] _IntNarrow_2_out;
/*mux_wire*/ logic _cur_start_chunk_addr_update;
/*mux_wire*/ logic[59:0] _cur_start_chunk_addr_new;
/*mux_wire*/ logic[32:0] next_num_chunks_left;
wire[8:0] _53;
assign _53 = next_arlen + 1'd1;
wire signed[33:0] _54;
assign _54 = __num_chunks_left_old_D0 - _53;
/*mux_wire*/ logic signed[33:0] _IntNarrow_3_in;
wire[32:0] _IntNarrow_3_out;
/*mux_wire*/ logic _num_chunks_left_update;
/*mux_wire*/ logic[32:0] _num_chunks_left_new;
/*mux_wire*/ logic _BoolToInt_i;
wire[0:0] _BoolToInt_o;
wire signed[12:0] _64;
assign _64 = num_in_flight - _BoolToInt_o;
wire _66;
assign _66 = !arvalid;
wire _68;
assign _68 = _66 & may_next_arvalid;
wire[8:0] _71;
assign _71 = next_arlen + 1'd1;
/*mux_wire*/ logic _Ternary_cond;
/*mux_wire*/ logic[8:0] _Ternary_a;
/*mux_wire*/ logic[8:0] _Ternary_b;
wire[8:0] _Ternary_o;
wire signed[12:0] _73;
assign _73 = _64 + $signed({1'b0, _Ternary_o});
/*mux_wire*/ logic signed[12:0] _IntNarrow_4_in;
wire[11:0] _IntNarrow_4_out;
/*state*/ logic[2:0] final_chunk_align;
/*state*/ logic[1:0] cur_chunk_align;
/*mux_wire*/ logic[31:0] elements_2[3:0];
wire[31:0] _75;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _75[_g0] = rdata[_g0];
end
endgenerate
wire[31:0] _76;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _76[_g0] = rdata[32 + _g0];
end
endgenerate
wire[31:0] _77;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _77[_g0] = rdata[64 + _g0];
end
endgenerate
wire[31:0] _78;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _78[_g0] = rdata[96 + _g0];
end
endgenerate
/*mux_wire*/ logic[2:0] num_chunk_elements;
/*mux_wire*/ logic is_last;
wire _81;
assign _81 = num_in_flight == 1'd1;
wire _83;
assign _83 = _81 & last_burst_in_flight;
wire signed[3:0] _87;
assign _87 = final_chunk_align - cur_chunk_align;
/*mux_wire*/ logic signed[3:0] _IntNarrow_5_in;
wire[2:0] _IntNarrow_5_out;
wire[2:0] _89;
assign _89 = 3'd4 - cur_chunk_align;
wire _97;
assign _97 = !chunks_are_left;
/*latency*/ logic __97_D0; always_ff @(posedge aclk) begin __97_D0 <= _97; end
wire _99;
assign _99 = __97_D0 & _num_chunks_left_may_update;
wire _101;
assign _101 = _99 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic[59:0] chunk_addr;
/*latency*/ logic[59:0] _chunk_addr_D1; always_ff @(posedge aclk) begin _chunk_addr_D1 <= chunk_addr; end
/*mux_wire*/ logic[1:0] element_in_chunk_align;
wire[61:0] _103;
assign _103 = start_addr / 3'd4;
/*mux_wire*/ logic[61:0] _BitwiseIntSplit_2_v;
wire[59:0] _BitwiseIntSplit_2_upper;
wire[1:0] _BitwiseIntSplit_2_lower;
/*mux_wire*/ logic[32:0] chunk_count_bits;
/*mux_wire*/ logic[1:0] final_alignment;
wire[34:0] _106;
assign _106 = count + element_in_chunk_align;
/*mux_wire*/ logic[34:0] _BitwiseIntSplit_3_v;
wire[32:0] _BitwiseIntSplit_3_upper;
wire[1:0] _BitwiseIntSplit_3_lower;
/*mux_wire*/ logic[32:0] num_chunks;
/*mux_wire*/ logic is_no_chunks;
wire _109;
assign _109 = chunk_count_bits == 1'd0;
wire _115;
assign _115 = final_alignment != 1'd0;
/*mux_wire*/ logic _BoolToInt_2_i;
wire[0:0] _BoolToInt_2_o;
wire[32:0] _116;
assign _116 = chunk_count_bits + _BoolToInt_2_o;
wire _122;
assign _122 = !is_no_chunks;
wire _125;
assign _125 = final_alignment == 1'd0;
wire _126;
assign _126 = _122 & _125;
/*mux_wire*/ logic _BoolToInt_3_i;
wire[0:0] _BoolToInt_3_o;
/*mux_wire*/ logic[0:0] _BitwiseIntConcat_3_upper;
/*mux_wire*/ logic[1:0] _BitwiseIntConcat_3_lower;
wire[2:0] _BitwiseIntConcat_3_v;
wire _130;
assign _130 = !aresetn;
/*mux_wire*/ logic _cur_start_chunk_addr_rst;
wire _132;
assign _132 = !aresetn;
/*mux_wire*/ logic _num_chunks_left_rst;
wire _134;
assign _134 = !aresetn;
SlowState_T_type_int_FROM_0_TO_1152921504606846976_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1 cur_start_chunk_addr(
	.clk(aclk),
	.rst(_cur_start_chunk_addr_rst),
	.old(_cur_start_chunk_addr_old),
	.may_update(_cur_start_chunk_addr_may_update),
	.update(_cur_start_chunk_addr_update),
	.new_1(_cur_start_chunk_addr_new)
);
SlowState_T_type_int_FROM_0_TO_4294967299_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0 num_chunks_left(
	.clk(aclk),
	.rst(_num_chunks_left_rst),
	.old(_num_chunks_left_old),
	.may_update(_num_chunks_left_may_update),
	.update(_num_chunks_left_update),
	.new_1(_num_chunks_left_new)
);
BitwiseIntConcat_UPPER_TO_1152921504606846976_LOWER_BITS_4 BitwiseIntConcat(
	.clk(aclk),
	.upper(_BitwiseIntConcat_upper),
	.lower(_BitwiseIntConcat_lower),
	.v(_BitwiseIntConcat_v)
);
BitwiseIntSplit_TO_1152921504606846976_LOWER_BITS_8 BitwiseIntSplit(
	.clk(aclk),
	.v(_BitwiseIntSplit_v),
	.upper(_BitwiseIntSplit_upper),
	.lower(_BitwiseIntSplit_lower)
);
IntNarrow_FROM_I_0_TO_I_4294967299_FROM_1_TO_257 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
LatencyOffset_T_type_bool_OFFSET_384 LatencyOffset(
	.clk(aclk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
BitwiseIntConcat_UPPER_TO_4503599627370497_LOWER_BITS_8 BitwiseIntConcat_2(
	.clk(aclk),
	.upper(_BitwiseIntConcat_2_upper),
	.lower(_BitwiseIntConcat_2_lower),
	.v(_BitwiseIntConcat_2_v)
);
IntNarrow_FROM_I_0_TO_I_1152921504606847232_FROM_0_TO_1152921504606846976 IntNarrow_2(
	.clk(aclk),
	.in(_IntNarrow_2_in),
	.out(_IntNarrow_2_out)
);
IntNarrow_FROM_I_256_TO_I_4294967298_FROM_0_TO_4294967299 IntNarrow_3(
	.clk(aclk),
	.in(_IntNarrow_3_in),
	.out(_IntNarrow_3_out)
);
BoolToInt BoolToInt(
	.clk(aclk),
	.i(_BoolToInt_i),
	.o(_BoolToInt_o)
);
Ternary_T_type_int_FROM_0_TO_257 Ternary(
	.clk(aclk),
	.cond(_Ternary_cond),
	.a(_Ternary_a),
	.b(_Ternary_b),
	.o(_Ternary_o)
);
IntNarrow_FROM_I_1_TO_I_3640_FROM_0_TO_3384 IntNarrow_4(
	.clk(aclk),
	.in(_IntNarrow_4_in),
	.out(_IntNarrow_4_out)
);
IntNarrow_FROM_I_3_TO_I_8_FROM_0_TO_5 IntNarrow_5(
	.clk(aclk),
	.in(_IntNarrow_5_in),
	.out(_IntNarrow_5_out)
);
BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_2 BitwiseIntSplit_2(
	.clk(aclk),
	.v(_BitwiseIntSplit_2_v),
	.upper(_BitwiseIntSplit_2_upper),
	.lower(_BitwiseIntSplit_2_lower)
);
BitwiseIntSplit_TO_17179869187_LOWER_BITS_2 BitwiseIntSplit_3(
	.clk(aclk),
	.v(_BitwiseIntSplit_3_v),
	.upper(_BitwiseIntSplit_3_upper),
	.lower(_BitwiseIntSplit_3_lower)
);
BoolToInt BoolToInt_2(
	.clk(aclk),
	.i(_BoolToInt_2_i),
	.o(_BoolToInt_2_o)
);
BoolToInt BoolToInt_3(
	.clk(aclk),
	.i(_BoolToInt_3_i),
	.o(_BoolToInt_3_o)
);
BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_2 BitwiseIntConcat_3(
	.clk(aclk),
	.upper(_BitwiseIntConcat_3_upper),
	.lower(_BitwiseIntConcat_3_lower),
	.v(_BitwiseIntConcat_3_v)
);
always_ff @(posedge aclk) begin // state arvalid
	if(arvalid) if(arready) arvalid <= 1'b0;
	if(!arvalid) if(may_next_arvalid) arvalid <= 1'b1;
	if(_134) arvalid <= 1'b0;
end
always_ff @(posedge aclk) begin // state araddr
	if(!arvalid) if(may_next_arvalid) araddr <= _next_araddr_D0;
end
always_ff @(posedge aclk) begin // state arlen
	if(!arvalid) if(may_next_arvalid) arlen <= next_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = 3'd4;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _1;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _2;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _3;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = 1'd0;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = 1'd0;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rresp = 2'bxx;
	_rresp = rresp;
end
always_comb begin // combinatorial _rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rlast = 1'bx;
	_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_rlast = _rlast;
end
always_comb begin // combinatorial element_packet_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_packet_valid = 1'bx;
	element_packet_valid = 1'b0;
	if(rvalid) element_packet_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	element_packet_valid = element_packet_valid;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
if(rvalid) elements[_v0] = elements_2[_v0];
end
end
always_comb begin // combinatorial chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_offset = 2'dx;
	if(rvalid) chunk_offset = cur_chunk_align;
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 3'dx;
	if(rvalid) chunk_length = num_chunk_elements;
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(rvalid) last = is_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state num_in_flight
	num_in_flight <= _IntNarrow_4_out;
	if(_134) num_in_flight <= 1'd0;
end
always_ff @(posedge aclk) begin // state last_burst_in_flight
	if(!arvalid) if(may_next_arvalid) last_burst_in_flight <= _next_last_burst_in_flight_D0;
end
always_comb begin // combinatorial next_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_araddr = 64'dx;
	next_araddr = _BitwiseIntConcat_v;
end
always_comb begin // combinatorial _BitwiseIntConcat_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_upper = 60'dx;
	_BitwiseIntConcat_upper = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial _BitwiseIntConcat_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_lower = 4'dx;
	_BitwiseIntConcat_lower = 1'd0;
end
always_comb begin // combinatorial next_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_arlen = 8'dx;
	if(_chunks_are_left_D0) if(__23_D0) next_arlen = __26_D0;
	if(_chunks_are_left_D0) if(!__23_D0) next_arlen = _max_chunks_in_this_burst_D0;
end
always_comb begin // combinatorial next_last_burst_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_last_burst_in_flight = 1'bx;
	next_last_burst_in_flight = 1'b0;
	if(chunks_are_left) if(_23) next_last_burst_in_flight = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	next_last_burst_in_flight = next_last_burst_in_flight;
end
always_comb begin // combinatorial cur_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_burst_addr = 52'dx;
	cur_burst_addr = _BitwiseIntSplit_upper;
end
always_comb begin // combinatorial cur_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_align = 8'dx;
	cur_align = _BitwiseIntSplit_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_v = 60'dx;
	_BitwiseIntSplit_v = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial chunks_are_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunks_are_left = 1'bx;
	chunks_are_left = __14_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunks_are_left = chunks_are_left;
end
always_comb begin // combinatorial max_chunks_in_this_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	max_chunks_in_this_burst = 8'dx;
	if(chunks_are_left) max_chunks_in_this_burst = _18;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 33'dx;
	if(chunks_are_left) if(_23) _IntNarrow_in = __num_chunks_left_old_N1;
end
always_comb begin // combinatorial may_next_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_next_arvalid = 1'bx;
	may_next_arvalid = _39;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_next_arvalid = may_next_arvalid;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial next_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_burst_addr = 53'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) next_burst_addr = __45_D1;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_upper = 53'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_upper = next_burst_addr;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_lower = 8'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_lower = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_2_in = 61'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _IntNarrow_2_in = _BitwiseIntConcat_2_v;
end
always_comb begin // combinatorial _cur_start_chunk_addr_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_update = 1'bx;
	_cur_start_chunk_addr_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _cur_start_chunk_addr_update = 1'b1;
	if(request_new_burst) _cur_start_chunk_addr_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_update = _cur_start_chunk_addr_update;
end
always_comb begin // combinatorial _cur_start_chunk_addr_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_new = 60'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _cur_start_chunk_addr_new = _IntNarrow_2_out;
	if(_request_new_burst_D1) _cur_start_chunk_addr_new = _chunk_addr_D1;
end
always_comb begin // combinatorial next_num_chunks_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_num_chunks_left = 33'dx;
	if(!arvalid) if(may_next_arvalid) next_num_chunks_left = _IntNarrow_3_out;
end
always_comb begin // combinatorial _IntNarrow_3_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_3_in = 34'sdx;
	if(!arvalid) if(may_next_arvalid) _IntNarrow_3_in = _54;
end
always_comb begin // combinatorial _num_chunks_left_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_update = 1'bx;
	_num_chunks_left_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_update = 1'b1;
	if(request_new_burst) _num_chunks_left_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_update = _num_chunks_left_update;
end
always_comb begin // combinatorial _num_chunks_left_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_new = 33'dx;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_new = next_num_chunks_left;
	if(request_new_burst) _num_chunks_left_new = num_chunks;
end
always_comb begin // combinatorial _BoolToInt_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_i = 1'bx;
	_BoolToInt_i = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_i = _BoolToInt_i;
end
always_comb begin // combinatorial _Ternary_cond
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_cond = 1'bx;
	_Ternary_cond = _68;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Ternary_cond = _Ternary_cond;
end
always_comb begin // combinatorial _Ternary_a
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_a = 9'dx;
	_Ternary_a = _71;
end
always_comb begin // combinatorial _Ternary_b
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_b = 9'dx;
	_Ternary_b = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_4_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_4_in = 13'sdx;
	_IntNarrow_4_in = _73;
end
always_ff @(posedge aclk) begin // state final_chunk_align
	if(request_new_burst) final_chunk_align <= _BitwiseIntConcat_3_v;
end
always_ff @(posedge aclk) begin // state cur_chunk_align
	if(rvalid) cur_chunk_align <= 1'd0;
	if(request_new_burst) cur_chunk_align <= element_in_chunk_align;
end
always_comb begin // combinatorial elements_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_2 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	if(rvalid) elements_2[0] = _75;
	if(rvalid) elements_2[1] = _76;
	if(rvalid) elements_2[2] = _77;
	if(rvalid) elements_2[3] = _78;
end
always_comb begin // combinatorial num_chunk_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunk_elements = 3'dx;
	if(rvalid) if(is_last) num_chunk_elements = _IntNarrow_5_out;
	if(rvalid) if(!is_last) num_chunk_elements = _89;
end
always_comb begin // combinatorial is_last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_last = 1'bx;
	if(rvalid) is_last = _83;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_last = is_last;
end
always_comb begin // combinatorial _IntNarrow_5_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_5_in = 4'sdx;
	if(rvalid) if(is_last) _IntNarrow_5_in = _87;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _101;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial chunk_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_addr = 60'dx;
	if(request_new_burst) chunk_addr = _BitwiseIntSplit_2_upper;
end
always_comb begin // combinatorial element_in_chunk_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_in_chunk_align = 2'dx;
	if(request_new_burst) element_in_chunk_align = _BitwiseIntSplit_2_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_2_v = 62'dx;
	if(request_new_burst) _BitwiseIntSplit_2_v = _103;
end
always_comb begin // combinatorial chunk_count_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_count_bits = 33'dx;
	if(request_new_burst) chunk_count_bits = _BitwiseIntSplit_3_upper;
end
always_comb begin // combinatorial final_alignment
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	final_alignment = 2'dx;
	if(request_new_burst) final_alignment = _BitwiseIntSplit_3_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_3_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_3_v = 35'dx;
	if(request_new_burst) _BitwiseIntSplit_3_v = _106;
end
always_comb begin // combinatorial num_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunks = 33'dx;
	if(request_new_burst) if(is_no_chunks) num_chunks = 1'd1;
	if(request_new_burst) if(!is_no_chunks) num_chunks = _116;
end
always_comb begin // combinatorial is_no_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_no_chunks = 1'bx;
	if(request_new_burst) is_no_chunks = _109;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_no_chunks = is_no_chunks;
end
always_comb begin // combinatorial _BoolToInt_2_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_2_i = 1'bx;
	if(request_new_burst) if(!is_no_chunks) _BoolToInt_2_i = _115;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_2_i = _BoolToInt_2_i;
end
always_comb begin // combinatorial _BoolToInt_3_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_3_i = 1'bx;
	if(request_new_burst) _BoolToInt_3_i = _126;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_3_i = _BoolToInt_3_i;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_upper = 1'dx;
	if(request_new_burst) _BitwiseIntConcat_3_upper = _BoolToInt_3_o;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BitwiseIntConcat_3_upper = _BitwiseIntConcat_3_upper;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_lower = 2'dx;
	if(request_new_burst) _BitwiseIntConcat_3_lower = final_alignment;
end
always_comb begin // combinatorial _cur_start_chunk_addr_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_rst = 1'bx;
	_cur_start_chunk_addr_rst = _130;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_rst = _cur_start_chunk_addr_rst;
end
always_comb begin // combinatorial _num_chunks_left_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_rst = 1'bx;
	_num_chunks_left_rst = _132;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_rst = _num_chunks_left_rst;
end
endmodule

// BitwiseIntSplit #(TO: 17179869187, LOWER_BITS: 2)
module BitwiseIntSplit_TO_17179869187_LOWER_BITS_2(
	input clk,
	input wire[34:0] v,
	output /*mux_wire*/ logic[32:0] upper,
	output /*mux_wire*/ logic[1:0] lower
);

genvar _g0;
/*mux_wire*/ logic[34:0] v_bits;
/*mux_wire*/ logic[34:0] _UIntToBits_value;
wire[34:0] _UIntToBits_bits;
wire[1:0] _2;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[1:0] _BitsToUInt_bits;
wire[1:0] _BitsToUInt_value;
wire[32:0] _3;
generate
for(_g0 = 0; _g0 < 33; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[2 + _g0];
end
endgenerate
/*mux_wire*/ logic[32:0] _FromBits_bits;
wire[32:0] _FromBits_value;
UIntToBits_NUM_BITS_35 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_2 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_4294967297 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 33'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 2'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 35'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 35'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 2'bxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// UIntToBits #(NUM_BITS: 35)
module UIntToBits_NUM_BITS_35(
	input clk,
	input wire[34:0] value,
	output /*mux_wire*/ logic[34:0] bits
);

	assign bits = value;
endmodule

// BitwiseIntSplit #(TO: 4611686018427387904, LOWER_BITS: 2)
module BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_2(
	input clk,
	input wire[61:0] v,
	output /*mux_wire*/ logic[59:0] upper,
	output /*mux_wire*/ logic[1:0] lower
);

genvar _g0;
/*mux_wire*/ logic[61:0] v_bits;
/*mux_wire*/ logic[61:0] _UIntToBits_value;
wire[61:0] _UIntToBits_bits;
wire[1:0] _2;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[1:0] _BitsToUInt_bits;
wire[1:0] _BitsToUInt_value;
wire[59:0] _3;
generate
for(_g0 = 0; _g0 < 60; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[2 + _g0];
end
endgenerate
/*mux_wire*/ logic[59:0] _FromBits_bits;
wire[59:0] _FromBits_value;
UIntToBits_NUM_BITS_62 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_2 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_1152921504606846976 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 60'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 2'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 62'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 62'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 2'bxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 60'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 1152921504606846976))
module FromBits_T_type_int_FROM_0_TO_1152921504606846976(
	input clk,
	input wire[59:0] bits,
	output /*mux_wire*/ logic[59:0] value
);

assign value = bits;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 1152921504606847232, FROM: 0, TO: 1152921504606846976)
module IntNarrow_FROM_I_0_TO_I_1152921504606847232_FROM_0_TO_1152921504606846976(
	input clk,
	input wire[60:0] in,
	output /*mux_wire*/ logic[59:0] out
);

	assign out = in;
endmodule

// BitwiseIntConcat #(UPPER_TO: 4503599627370497, LOWER_BITS: 8)
module BitwiseIntConcat_UPPER_TO_4503599627370497_LOWER_BITS_8(
	input clk,
	input wire[52:0] upper,
	input wire[7:0] lower,
	output /*mux_wire*/ logic[60:0] v
);

/*mux_wire*/ logic[60:0] v_bits;
/*mux_wire*/ logic[7:0] _UIntToBits_value;
wire[7:0] _UIntToBits_bits;
/*mux_wire*/ logic[52:0] _UIntToBits_2_value;
wire[52:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[60:0] _FromBits_bits;
wire[60:0] _FromBits_value;
UIntToBits_NUM_BITS_8 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_53 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_1152921504606847232 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 61'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 61'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 53; _v0 = _v0 + 1) begin
v_bits[8 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 8'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 53'dx;
	_UIntToBits_2_value = upper;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 61'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 1152921504606847232))
module FromBits_T_type_int_FROM_0_TO_1152921504606847232(
	input clk,
	input wire[60:0] bits,
	output /*mux_wire*/ logic[60:0] value
);

assign value = bits;
endmodule

// BitwiseIntSplit #(TO: 1152921504606846976, LOWER_BITS: 8)
module BitwiseIntSplit_TO_1152921504606846976_LOWER_BITS_8(
	input clk,
	input wire[59:0] v,
	output /*mux_wire*/ logic[51:0] upper,
	output /*mux_wire*/ logic[7:0] lower
);

genvar _g0;
/*mux_wire*/ logic[59:0] v_bits;
/*mux_wire*/ logic[59:0] _UIntToBits_value;
wire[59:0] _UIntToBits_bits;
wire[7:0] _2;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[7:0] _BitsToUInt_bits;
wire[7:0] _BitsToUInt_value;
wire[51:0] _3;
generate
for(_g0 = 0; _g0 < 52; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[8 + _g0];
end
endgenerate
/*mux_wire*/ logic[51:0] _FromBits_bits;
wire[51:0] _FromBits_value;
UIntToBits_NUM_BITS_60 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_8 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_4503599627370496 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 52'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 8'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 60'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 60'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 8'bxxxxxxxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 52'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// BitwiseIntConcat #(UPPER_TO: 1152921504606846976, LOWER_BITS: 4)
module BitwiseIntConcat_UPPER_TO_1152921504606846976_LOWER_BITS_4(
	input clk,
	input wire[59:0] upper,
	input wire[3:0] lower,
	output /*mux_wire*/ logic[63:0] v
);

/*mux_wire*/ logic[63:0] v_bits;
/*mux_wire*/ logic[3:0] _UIntToBits_value;
wire[3:0] _UIntToBits_bits;
/*mux_wire*/ logic[59:0] _UIntToBits_2_value;
wire[59:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[63:0] _FromBits_bits;
wire[63:0] _FromBits_value;
UIntToBits_NUM_BITS_4 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_60 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_18446744073709551616 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 64'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 60; _v0 = _v0 + 1) begin
v_bits[4 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 4'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 60'dx;
	_UIntToBits_2_value = upper;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// UIntToBits #(NUM_BITS: 60)
module UIntToBits_NUM_BITS_60(
	input clk,
	input wire[59:0] value,
	output /*mux_wire*/ logic[59:0] bits
);

	assign bits = value;
endmodule

// SlowState #(T: type int #(FROM: 0, TO: 1152921504606846976), RESET_TO: 0, OLD_DELAY: 1, NEW_DELAY: 1)
module SlowState_T_type_int_FROM_0_TO_1152921504606846976_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1(
	input clk,
	input wire rst,
	output /*state*/ logic[59:0] old,
	output /*mux_wire*/ logic may_update,
	input wire update,
	input wire[59:0] new_1
);

/*latency*/ logic _update_D1; always_ff @(posedge clk) begin _update_D1 <= update; end
genvar _g0;
/*mux_wire*/ logic _cross_rst_in;
/*mux_wire*/ logic[59:0] new_s;
/*mux_wire*/ logic update_s;
/*mux_wire*/ logic update_old;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
/*latency*/ logic __LatencyOffset_out_N1; always_ff @(posedge clk) begin __LatencyOffset_out_N1 <= _LatencyOffset_out; end
/*mux_wire*/ logic[59:0] new_old;
/*mux_wire*/ logic[59:0] _LatencyOffset_2_in;
wire[59:0] _LatencyOffset_2_out;
wire _cross_rst_out;
/*latency*/ logic __cross_rst_out_D0; always_ff @(posedge clk) begin __cross_rst_out_D0 <= _cross_rst_out; end
/*state*/ logic[1:0] cooldown;
wire _8 = cooldown[0];
wire _11;
assign _11 = update_s | __cross_rst_out_D0;
/*mux_wire*/ logic _Repeat_v;
wire[1:0] _Repeat_result;
wire[0:0] _12;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _12[_g0] = cooldown[1 + _g0];
end
endgenerate
CrossDomain_T_type_bool cross_rst(
	.in_clk(clk),
	.in(_cross_rst_in),
	.out(_cross_rst_out)
);
LatencyOffset_T_type_bool_OFFSET_2 LatencyOffset(
	.clk(clk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
LatencyOffset_T_type_int_FROM_0_TO_1152921504606846976_OFFSET_2 LatencyOffset_2(
	.clk(clk),
	.in(_LatencyOffset_2_in),
	.out(_LatencyOffset_2_out)
);
Repeat_T_type_bool_SIZE_2 Repeat(
	.clk(clk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
always_comb begin // combinatorial _cross_rst_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_rst_in = 1'bx;
	_cross_rst_in = rst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_rst_in = _cross_rst_in;
end
always_ff @(posedge clk) begin // state old
	if(_cross_rst_out) old <= 60'd0;
	if(!_cross_rst_out) if(update_old) old <= new_old;
end
always_comb begin // combinatorial new_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_s = 60'dx;
	if(_update_D1) new_s = new_1;
end
always_comb begin // combinatorial update_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_s = 1'bx;
	if(update) update_s = 1'b1;
	if(!update) update_s = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_s = update_s;
end
always_comb begin // combinatorial update_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_old = 1'bx;
	update_old = __LatencyOffset_out_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_old = update_old;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = update_s;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial new_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_old = 60'dx;
	new_old = _LatencyOffset_2_out;
end
always_comb begin // combinatorial _LatencyOffset_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_2_in = 60'dx;
	_LatencyOffset_2_in = new_s;
end
always_comb begin // combinatorial may_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_update = 1'bx;
	may_update = _8;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_update = may_update;
end
always_ff @(posedge clk) begin // state cooldown
	if(_11) cooldown <= _Repeat_result;
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(!_11) cooldown[_v0] <= _12[_v0];
end
	if(!_11) cooldown[1] <= 1'b1;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	if(_11) _Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
endmodule

// LatencyOffset #(T: type int #(FROM: 0, TO: 1152921504606846976), OFFSET: -2)
module LatencyOffset_T_type_int_FROM_0_TO_1152921504606846976_OFFSET_2(
	input clk,
	input wire[59:0] in,
	output /*mux_wire*/ logic[59:0] out
);

	assign out = in;
endmodule

// benchmark_burst_read #(AXI_WIDTH: 64)
module benchmark_burst_read_AXI_WIDTH_64(
	input aclk,
	input wire aresetn,
	input wire[11:0] s_axi_control_awaddr,
	input wire s_axi_control_awvalid,
	output /*mux_wire*/ logic s_axi_control_awready,
	input wire[31:0] s_axi_control_wdata,
	input wire[3:0] s_axi_control_wstrb,
	input wire s_axi_control_wvalid,
	output /*mux_wire*/ logic s_axi_control_wready,
	output /*mux_wire*/ logic[1:0] s_axi_control_bresp,
	output /*mux_wire*/ logic s_axi_control_bvalid,
	input wire s_axi_control_bready,
	input wire[11:0] s_axi_control_araddr,
	input wire s_axi_control_arvalid,
	output /*mux_wire*/ logic s_axi_control_arready,
	output /*mux_wire*/ logic[31:0] s_axi_control_rdata,
	output /*mux_wire*/ logic[1:0] s_axi_control_rresp,
	output /*mux_wire*/ logic s_axi_control_rvalid,
	input wire s_axi_control_rready,
	output /*mux_wire*/ logic m_axi_awvalid,
	input wire m_axi_awready,
	output /*mux_wire*/ logic[63:0] m_axi_awaddr,
	output /*mux_wire*/ logic[7:0] m_axi_awlen,
	output /*mux_wire*/ logic[1:0] m_axi_awburst,
	output /*mux_wire*/ logic[3:0] m_axi_awcache,
	output /*mux_wire*/ logic m_axi_wvalid,
	input wire m_axi_wready,
	output /*mux_wire*/ logic[63:0] m_axi_wdata,
	output /*mux_wire*/ logic[7:0] m_axi_wstrb,
	output /*mux_wire*/ logic m_axi_wlast,
	input wire m_axi_bvalid,
	output /*mux_wire*/ logic m_axi_bready,
	input wire[1:0] m_axi_bresp,
	output /*mux_wire*/ logic m_axi_arvalid,
	input wire m_axi_arready,
	output /*mux_wire*/ logic[63:0] m_axi_araddr,
	output /*mux_wire*/ logic[7:0] m_axi_arlen,
	output /*mux_wire*/ logic[2:0] m_axi_arsize,
	output /*mux_wire*/ logic[1:0] m_axi_arburst,
	input wire m_axi_rvalid,
	output /*mux_wire*/ logic m_axi_rready,
	input wire[63:0] m_axi_rdata,
	input wire[1:0] m_axi_rresp,
	input wire m_axi_rlast,
	output /*mux_wire*/ logic[2:0] m_axi_arprot,
	output /*mux_wire*/ logic[3:0] m_axi_arcache,
	output /*mux_wire*/ logic[3:0] m_axi_arqos,
	output /*mux_wire*/ logic m_axi_arlock,
	output /*mux_wire*/ logic[3:0] m_axi_arregion
);

genvar _g0;
/*mux_wire*/ logic _ctrl_aresetn;
wire _ctrl_awready;
wire _ctrl_wready;
wire[1:0] _ctrl_bresp;
wire _ctrl_bvalid;
wire _ctrl_arready;
wire[31:0] _ctrl_rdata;
wire[1:0] _ctrl_rresp;
wire _ctrl_rvalid;
/*mux_wire*/ logic[11:0] _ctrl_awaddr;
/*mux_wire*/ logic _ctrl_awvalid;
/*mux_wire*/ logic[31:0] _ctrl_wdata;
/*mux_wire*/ logic[3:0] _ctrl_wstrb;
/*mux_wire*/ logic _ctrl_wvalid;
/*mux_wire*/ logic _ctrl_bready;
/*mux_wire*/ logic[11:0] _ctrl_araddr;
/*mux_wire*/ logic _ctrl_arvalid;
/*mux_wire*/ logic _ctrl_rready;
/*mux_wire*/ logic _reader_aresetn;
/*mux_wire*/ logic _writer_aresetn;
wire _writer_awvalid;
wire[63:0] _writer_awaddr;
wire[7:0] _writer_awlen;
wire[1:0] _writer_awburst;
wire[3:0] _writer_awcache;
wire _writer_wvalid;
wire[63:0] _writer_wdata;
wire[7:0] _writer_wstrb;
wire _writer_wlast;
wire _writer_bready;
/*mux_wire*/ logic _writer_awready;
/*mux_wire*/ logic _writer_wready;
/*mux_wire*/ logic _writer_bvalid;
/*mux_wire*/ logic[1:0] _writer_bresp;
wire _reader_arvalid;
wire[63:0] _reader_araddr;
wire[7:0] _reader_arlen;
wire[2:0] _reader_arsize;
wire[1:0] _reader_arburst;
wire _reader_rready;
/*mux_wire*/ logic _reader_arready;
/*mux_wire*/ logic _reader_rvalid;
/*mux_wire*/ logic[63:0] _reader_rdata;
/*mux_wire*/ logic[1:0] _reader_rresp;
/*mux_wire*/ logic _reader_rlast;
/*mux_wire*/ logic[63:0] addr_a_bits;
wire[31:0] _ctrl_input_regs[3:0];
wire[31:0] _46 = _ctrl_input_regs[0];
wire[31:0] _47 = _ctrl_input_regs[1];
/*mux_wire*/ logic[63:0] start_addr;
/*mux_wire*/ logic[63:0] _BitsToUInt_bits;
wire[63:0] _BitsToUInt_value;
/*mux_wire*/ logic[31:0] num_to_transfer;
wire[31:0] _49 = _ctrl_input_regs[2];
/*mux_wire*/ logic[31:0] _BitsToUInt_2_bits;
wire[31:0] _BitsToUInt_2_value;
/*mux_wire*/ logic[31:0] _IntNarrow_in;
wire[31:0] _IntNarrow_out;
/*mux_wire*/ logic[31:0] config_bits;
wire[31:0] _50 = _ctrl_input_regs[3];
wire[2:0] _51;
generate
for(_g0 = 0; _g0 < 3; _g0 = _g0 + 1) begin
assign _51[_g0] = config_bits[5 + _g0];
end
endgenerate
wire[3:0] _52;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _52[_g0] = config_bits[8 + _g0];
end
endgenerate
wire[3:0] _53;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _53[_g0] = config_bits[12 + _g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_3_bits;
wire[3:0] _BitsToUInt_3_value;
wire _54 = config_bits[16];
wire[3:0] _55;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _55[_g0] = config_bits[17 + _g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_4_bits;
wire[3:0] _BitsToUInt_4_value;
wire[10:0] _56;
generate
for(_g0 = 0; _g0 < 11; _g0 = _g0 + 1) begin
assign _56[_g0] = config_bits[21 + _g0];
end
endgenerate
/*mux_wire*/ logic[10:0] _BitsToUInt_5_bits;
wire[10:0] _BitsToUInt_5_value;
/*mux_wire*/ logic[10:0] _reader_max_in_flight;
/*state*/ logic[63:0] cycles_since_reset;
wire[64:0] _59;
assign _59 = cycles_since_reset + 1'd1;
wire[63:0] _60;
assign _60 = _59; // == mod 18446744073709551616 (target is 64 bits wide)
/*mux_wire*/ logic[63:0] cycles_since_reset_bits;
/*mux_wire*/ logic[63:0] _UIntToBits_value;
wire[63:0] _UIntToBits_bits;
/*latency*/ logic[63:0] __UIntToBits_bits_D1; always_ff @(posedge aclk) begin __UIntToBits_bits_D1 <= _UIntToBits_bits; end
/*latency*/ logic[63:0] __UIntToBits_bits_D2; always_ff @(posedge aclk) begin __UIntToBits_bits_D2 <= __UIntToBits_bits_D1; end
/*latency*/ logic[63:0] __UIntToBits_bits_D3; always_ff @(posedge aclk) begin __UIntToBits_bits_D3 <= __UIntToBits_bits_D2; end
/*state*/ logic[63:0] cycles_since_reset_at_start;
/*state*/ logic running;
/*state*/ logic[31:0] num_cycles_running;
/*state*/ logic[31:0] hash;
wire _ctrl_start;
/*latency*/ logic __ctrl_start_D1; always_ff @(posedge aclk) begin __ctrl_start_D1 <= _ctrl_start; end
/*latency*/ logic __ctrl_start_D2; always_ff @(posedge aclk) begin __ctrl_start_D2 <= __ctrl_start_D1; end
/*latency*/ logic __ctrl_start_D3; always_ff @(posedge aclk) begin __ctrl_start_D3 <= __ctrl_start_D2; end
/*mux_wire*/ logic _reader_request_new_burst;
/*mux_wire*/ logic[63:0] _reader_start_addr;
/*mux_wire*/ logic[31:0] _reader_count;
localparam[31:0] _67 = 32'b00000000000000000000000000000000;
wire[32:0] _72;
assign _72 = num_cycles_running + 1'd1;
wire[31:0] _73;
assign _73 = _72; // == mod 4294967296 (target is 32 bits wide)
/*mux_wire*/ logic _reader_is_ready_to_receive_lots_of_data;
wire _reader_value_valid;
/*latency*/ logic __reader_value_valid_D1; always_ff @(posedge aclk) begin __reader_value_valid_D1 <= _reader_value_valid; end
/*latency*/ logic __reader_value_valid_D2; always_ff @(posedge aclk) begin __reader_value_valid_D2 <= __reader_value_valid_D1; end
/*latency*/ logic __reader_value_valid_D3; always_ff @(posedge aclk) begin __reader_value_valid_D3 <= __reader_value_valid_D2; end
wire[31:0] _reader_value[1:0];
wire _reader_last;
/*mux_wire*/ logic[31:0] value[1:0];
/*mux_wire*/ logic last;
/*latency*/ logic _last_D1; always_ff @(posedge aclk) begin _last_D1 <= last; end
/*latency*/ logic _last_D2; always_ff @(posedge aclk) begin _last_D2 <= _last_D1; end
/*latency*/ logic _last_D3; always_ff @(posedge aclk) begin _last_D3 <= _last_D2; end
/*mux_wire*/ logic[31:0] new_hash_contrib;
wire[1:0] _74;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _74[_g0] = value[_g0][0];
end
endgenerate
wire _75;
assign _75 = ^_74;
/*latency*/ logic __75_D1; always_ff @(posedge aclk) begin __75_D1 <= _75; end
/*latency*/ logic __75_D2; always_ff @(posedge aclk) begin __75_D2 <= __75_D1; end
wire[1:0] _76;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _76[_g0] = value[_g0][1];
end
endgenerate
wire _77;
assign _77 = ^_76;
/*latency*/ logic __77_D1; always_ff @(posedge aclk) begin __77_D1 <= _77; end
/*latency*/ logic __77_D2; always_ff @(posedge aclk) begin __77_D2 <= __77_D1; end
wire[1:0] _78;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _78[_g0] = value[_g0][2];
end
endgenerate
wire _79;
assign _79 = ^_78;
/*latency*/ logic __79_D1; always_ff @(posedge aclk) begin __79_D1 <= _79; end
/*latency*/ logic __79_D2; always_ff @(posedge aclk) begin __79_D2 <= __79_D1; end
wire[1:0] _80;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _80[_g0] = value[_g0][3];
end
endgenerate
wire _81;
assign _81 = ^_80;
/*latency*/ logic __81_D1; always_ff @(posedge aclk) begin __81_D1 <= _81; end
/*latency*/ logic __81_D2; always_ff @(posedge aclk) begin __81_D2 <= __81_D1; end
wire[1:0] _82;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _82[_g0] = value[_g0][4];
end
endgenerate
wire _83;
assign _83 = ^_82;
/*latency*/ logic __83_D1; always_ff @(posedge aclk) begin __83_D1 <= _83; end
/*latency*/ logic __83_D2; always_ff @(posedge aclk) begin __83_D2 <= __83_D1; end
wire[1:0] _84;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _84[_g0] = value[_g0][5];
end
endgenerate
wire _85;
assign _85 = ^_84;
/*latency*/ logic __85_D1; always_ff @(posedge aclk) begin __85_D1 <= _85; end
/*latency*/ logic __85_D2; always_ff @(posedge aclk) begin __85_D2 <= __85_D1; end
wire[1:0] _86;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _86[_g0] = value[_g0][6];
end
endgenerate
wire _87;
assign _87 = ^_86;
/*latency*/ logic __87_D1; always_ff @(posedge aclk) begin __87_D1 <= _87; end
/*latency*/ logic __87_D2; always_ff @(posedge aclk) begin __87_D2 <= __87_D1; end
wire[1:0] _88;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _88[_g0] = value[_g0][7];
end
endgenerate
wire _89;
assign _89 = ^_88;
/*latency*/ logic __89_D1; always_ff @(posedge aclk) begin __89_D1 <= _89; end
/*latency*/ logic __89_D2; always_ff @(posedge aclk) begin __89_D2 <= __89_D1; end
wire[1:0] _90;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _90[_g0] = value[_g0][8];
end
endgenerate
wire _91;
assign _91 = ^_90;
/*latency*/ logic __91_D1; always_ff @(posedge aclk) begin __91_D1 <= _91; end
/*latency*/ logic __91_D2; always_ff @(posedge aclk) begin __91_D2 <= __91_D1; end
wire[1:0] _92;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _92[_g0] = value[_g0][9];
end
endgenerate
wire _93;
assign _93 = ^_92;
/*latency*/ logic __93_D1; always_ff @(posedge aclk) begin __93_D1 <= _93; end
/*latency*/ logic __93_D2; always_ff @(posedge aclk) begin __93_D2 <= __93_D1; end
wire[1:0] _94;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _94[_g0] = value[_g0][10];
end
endgenerate
wire _95;
assign _95 = ^_94;
/*latency*/ logic __95_D1; always_ff @(posedge aclk) begin __95_D1 <= _95; end
/*latency*/ logic __95_D2; always_ff @(posedge aclk) begin __95_D2 <= __95_D1; end
wire[1:0] _96;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _96[_g0] = value[_g0][11];
end
endgenerate
wire _97;
assign _97 = ^_96;
/*latency*/ logic __97_D1; always_ff @(posedge aclk) begin __97_D1 <= _97; end
/*latency*/ logic __97_D2; always_ff @(posedge aclk) begin __97_D2 <= __97_D1; end
wire[1:0] _98;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _98[_g0] = value[_g0][12];
end
endgenerate
wire _99;
assign _99 = ^_98;
/*latency*/ logic __99_D1; always_ff @(posedge aclk) begin __99_D1 <= _99; end
/*latency*/ logic __99_D2; always_ff @(posedge aclk) begin __99_D2 <= __99_D1; end
wire[1:0] _100;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _100[_g0] = value[_g0][13];
end
endgenerate
wire _101;
assign _101 = ^_100;
/*latency*/ logic __101_D1; always_ff @(posedge aclk) begin __101_D1 <= _101; end
/*latency*/ logic __101_D2; always_ff @(posedge aclk) begin __101_D2 <= __101_D1; end
wire[1:0] _102;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _102[_g0] = value[_g0][14];
end
endgenerate
wire _103;
assign _103 = ^_102;
/*latency*/ logic __103_D1; always_ff @(posedge aclk) begin __103_D1 <= _103; end
/*latency*/ logic __103_D2; always_ff @(posedge aclk) begin __103_D2 <= __103_D1; end
wire[1:0] _104;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _104[_g0] = value[_g0][15];
end
endgenerate
wire _105;
assign _105 = ^_104;
/*latency*/ logic __105_D1; always_ff @(posedge aclk) begin __105_D1 <= _105; end
/*latency*/ logic __105_D2; always_ff @(posedge aclk) begin __105_D2 <= __105_D1; end
wire[1:0] _106;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _106[_g0] = value[_g0][16];
end
endgenerate
wire _107;
assign _107 = ^_106;
/*latency*/ logic __107_D1; always_ff @(posedge aclk) begin __107_D1 <= _107; end
/*latency*/ logic __107_D2; always_ff @(posedge aclk) begin __107_D2 <= __107_D1; end
wire[1:0] _108;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _108[_g0] = value[_g0][17];
end
endgenerate
wire _109;
assign _109 = ^_108;
/*latency*/ logic __109_D1; always_ff @(posedge aclk) begin __109_D1 <= _109; end
/*latency*/ logic __109_D2; always_ff @(posedge aclk) begin __109_D2 <= __109_D1; end
wire[1:0] _110;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _110[_g0] = value[_g0][18];
end
endgenerate
wire _111;
assign _111 = ^_110;
/*latency*/ logic __111_D1; always_ff @(posedge aclk) begin __111_D1 <= _111; end
/*latency*/ logic __111_D2; always_ff @(posedge aclk) begin __111_D2 <= __111_D1; end
wire[1:0] _112;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _112[_g0] = value[_g0][19];
end
endgenerate
wire _113;
assign _113 = ^_112;
/*latency*/ logic __113_D1; always_ff @(posedge aclk) begin __113_D1 <= _113; end
/*latency*/ logic __113_D2; always_ff @(posedge aclk) begin __113_D2 <= __113_D1; end
wire[1:0] _114;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _114[_g0] = value[_g0][20];
end
endgenerate
wire _115;
assign _115 = ^_114;
/*latency*/ logic __115_D1; always_ff @(posedge aclk) begin __115_D1 <= _115; end
/*latency*/ logic __115_D2; always_ff @(posedge aclk) begin __115_D2 <= __115_D1; end
wire[1:0] _116;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _116[_g0] = value[_g0][21];
end
endgenerate
wire _117;
assign _117 = ^_116;
/*latency*/ logic __117_D1; always_ff @(posedge aclk) begin __117_D1 <= _117; end
/*latency*/ logic __117_D2; always_ff @(posedge aclk) begin __117_D2 <= __117_D1; end
wire[1:0] _118;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _118[_g0] = value[_g0][22];
end
endgenerate
wire _119;
assign _119 = ^_118;
/*latency*/ logic __119_D1; always_ff @(posedge aclk) begin __119_D1 <= _119; end
/*latency*/ logic __119_D2; always_ff @(posedge aclk) begin __119_D2 <= __119_D1; end
wire[1:0] _120;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _120[_g0] = value[_g0][23];
end
endgenerate
wire _121;
assign _121 = ^_120;
/*latency*/ logic __121_D1; always_ff @(posedge aclk) begin __121_D1 <= _121; end
/*latency*/ logic __121_D2; always_ff @(posedge aclk) begin __121_D2 <= __121_D1; end
wire[1:0] _122;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _122[_g0] = value[_g0][24];
end
endgenerate
wire _123;
assign _123 = ^_122;
/*latency*/ logic __123_D1; always_ff @(posedge aclk) begin __123_D1 <= _123; end
/*latency*/ logic __123_D2; always_ff @(posedge aclk) begin __123_D2 <= __123_D1; end
wire[1:0] _124;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _124[_g0] = value[_g0][25];
end
endgenerate
wire _125;
assign _125 = ^_124;
/*latency*/ logic __125_D1; always_ff @(posedge aclk) begin __125_D1 <= _125; end
/*latency*/ logic __125_D2; always_ff @(posedge aclk) begin __125_D2 <= __125_D1; end
wire[1:0] _126;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _126[_g0] = value[_g0][26];
end
endgenerate
wire _127;
assign _127 = ^_126;
/*latency*/ logic __127_D1; always_ff @(posedge aclk) begin __127_D1 <= _127; end
/*latency*/ logic __127_D2; always_ff @(posedge aclk) begin __127_D2 <= __127_D1; end
wire[1:0] _128;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _128[_g0] = value[_g0][27];
end
endgenerate
wire _129;
assign _129 = ^_128;
/*latency*/ logic __129_D1; always_ff @(posedge aclk) begin __129_D1 <= _129; end
/*latency*/ logic __129_D2; always_ff @(posedge aclk) begin __129_D2 <= __129_D1; end
wire[1:0] _130;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _130[_g0] = value[_g0][28];
end
endgenerate
wire _131;
assign _131 = ^_130;
/*latency*/ logic __131_D1; always_ff @(posedge aclk) begin __131_D1 <= _131; end
/*latency*/ logic __131_D2; always_ff @(posedge aclk) begin __131_D2 <= __131_D1; end
wire[1:0] _132;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _132[_g0] = value[_g0][29];
end
endgenerate
wire _133;
assign _133 = ^_132;
/*latency*/ logic __133_D1; always_ff @(posedge aclk) begin __133_D1 <= _133; end
/*latency*/ logic __133_D2; always_ff @(posedge aclk) begin __133_D2 <= __133_D1; end
wire[1:0] _134;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _134[_g0] = value[_g0][30];
end
endgenerate
wire _135;
assign _135 = ^_134;
/*latency*/ logic __135_D1; always_ff @(posedge aclk) begin __135_D1 <= _135; end
/*latency*/ logic __135_D2; always_ff @(posedge aclk) begin __135_D2 <= __135_D1; end
wire[1:0] _136;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _136[_g0] = value[_g0][31];
end
endgenerate
wire _137;
assign _137 = ^_136;
/*latency*/ logic __137_D1; always_ff @(posedge aclk) begin __137_D1 <= _137; end
/*latency*/ logic __137_D2; always_ff @(posedge aclk) begin __137_D2 <= __137_D1; end
/*mux_wire*/ logic[31:0] new_hash;
/*latency*/ logic[31:0] _new_hash_D3; always_ff @(posedge aclk) begin _new_hash_D3 <= new_hash; end
wire[31:0] _140;
assign _140 = hash ^ new_hash_contrib;
/*mux_wire*/ logic[31:0] _UIntToBits_2_value;
wire[31:0] _UIntToBits_2_bits;
/*latency*/ logic[31:0] __UIntToBits_2_bits_D1; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D1 <= _UIntToBits_2_bits; end
/*latency*/ logic[31:0] __UIntToBits_2_bits_D2; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D2 <= __UIntToBits_2_bits_D1; end
/*latency*/ logic[31:0] __UIntToBits_2_bits_D3; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D3 <= __UIntToBits_2_bits_D2; end
wire[31:0] _144;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _144[_g0] = cycles_since_reset_at_start[_g0];
end
endgenerate
wire[31:0] _145;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _145[_g0] = cycles_since_reset_at_start[32 + _g0];
end
endgenerate
wire[31:0] _146;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _146[_g0] = cycles_since_reset_bits[_g0];
end
endgenerate
wire[31:0] _147;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _147[_g0] = cycles_since_reset_bits[32 + _g0];
end
endgenerate
wire[31:0] _148[5:0];
assign _148[0] = __UIntToBits_2_bits_D3;
assign _148[1] = _new_hash_D3;
assign _148[2] = _144;
assign _148[3] = _145;
assign _148[4] = _146;
assign _148[5] = _147;
/*mux_wire*/ logic _ctrl_finish;
/*mux_wire*/ logic[31:0] _ctrl_output_regs[5:0];
wire _153;
assign _153 = !aresetn;
/*latency*/ logic __153_D1; always_ff @(posedge aclk) begin __153_D1 <= _153; end
/*latency*/ logic __153_D2; always_ff @(posedge aclk) begin __153_D2 <= __153_D1; end
localparam[31:0] _155 = 32'b00000000000000000000000000000000;
axi_ctrl_slave_NUM_INPUT_REGS_4_NUM_OUTPUT_REGS_6_ADDR_WIDTH_12_AXI_WIDTH_32 ctrl(
	.aclk(aclk),
	.aresetn(_ctrl_aresetn),
	.awaddr(_ctrl_awaddr),
	.awvalid(_ctrl_awvalid),
	.awready(_ctrl_awready),
	.wdata(_ctrl_wdata),
	.wstrb(_ctrl_wstrb),
	.wvalid(_ctrl_wvalid),
	.wready(_ctrl_wready),
	.bresp(_ctrl_bresp),
	.bvalid(_ctrl_bvalid),
	.bready(_ctrl_bready),
	.araddr(_ctrl_araddr),
	.arvalid(_ctrl_arvalid),
	.arready(_ctrl_arready),
	.rdata(_ctrl_rdata),
	.rresp(_ctrl_rresp),
	.rvalid(_ctrl_rvalid),
	.rready(_ctrl_rready),
	.input_regs(_ctrl_input_regs),
	.start(_ctrl_start),
	.finish(_ctrl_finish),
	.output_regs(_ctrl_output_regs)
);
axi_realigning_burst_reader_T_type_bool_32_2_AXI_WIDTH_64_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616 reader(
	.aclk(aclk),
	.aresetn(_reader_aresetn),
	.arvalid(_reader_arvalid),
	.arready(_reader_arready),
	.araddr(_reader_araddr),
	.arlen(_reader_arlen),
	.arsize(_reader_arsize),
	.arburst(_reader_arburst),
	.arprot(),
	.arcache(),
	.arqos(),
	.arlock(),
	.arregion(),
	.rvalid(_reader_rvalid),
	.rready(_reader_rready),
	.rdata(_reader_rdata),
	.rresp(_reader_rresp),
	.rlast(_reader_rlast),
	.max_in_flight(_reader_max_in_flight),
	.may_request_new_burst(),
	.request_new_burst(_reader_request_new_burst),
	.start_addr(_reader_start_addr),
	.count(_reader_count),
	.is_ready_to_receive_lots_of_data(_reader_is_ready_to_receive_lots_of_data),
	.value_valid(_reader_value_valid),
	.value(_reader_value),
	.last(_reader_last)
);
axi_memory_writer_tie_off_AXI_WIDTH_64 writer(
	.aclk(aclk),
	.aresetn(_writer_aresetn),
	.awvalid(_writer_awvalid),
	.awready(_writer_awready),
	.awaddr(_writer_awaddr),
	.awlen(_writer_awlen),
	.awsize(),
	.awburst(_writer_awburst),
	.awprot(),
	.awcache(_writer_awcache),
	.awqos(),
	.awlock(),
	.awregion(),
	.wvalid(_writer_wvalid),
	.wready(_writer_wready),
	.wdata(_writer_wdata),
	.wstrb(_writer_wstrb),
	.wlast(_writer_wlast),
	.bvalid(_writer_bvalid),
	.bresp(_writer_bresp),
	.bready(_writer_bready)
);
BitsToUInt_NUM_BITS_64 BitsToUInt(
	.clk(aclk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
BitsToUInt_NUM_BITS_32 BitsToUInt_2(
	.clk(aclk),
	.bits(_BitsToUInt_2_bits),
	.value(_BitsToUInt_2_value)
);
IntNarrow_FROM_I_0_TO_I_4294967296_FROM_1_TO_4294967296 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
BitsToUInt_NUM_BITS_4 BitsToUInt_3(
	.clk(aclk),
	.bits(_BitsToUInt_3_bits),
	.value(_BitsToUInt_3_value)
);
BitsToUInt_NUM_BITS_4 BitsToUInt_4(
	.clk(aclk),
	.bits(_BitsToUInt_4_bits),
	.value(_BitsToUInt_4_value)
);
BitsToUInt_NUM_BITS_11 BitsToUInt_5(
	.clk(aclk),
	.bits(_BitsToUInt_5_bits),
	.value(_BitsToUInt_5_value)
);
UIntToBits_NUM_BITS_64 UIntToBits(
	.clk(aclk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_32 UIntToBits_2(
	.clk(aclk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
always_comb begin // combinatorial _ctrl_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_aresetn = 1'bx;
	_ctrl_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_aresetn = _ctrl_aresetn;
end
always_comb begin // combinatorial s_axi_control_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_awready = 1'bx;
	s_axi_control_awready = _ctrl_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_awready = s_axi_control_awready;
end
always_comb begin // combinatorial s_axi_control_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_wready = 1'bx;
	s_axi_control_wready = _ctrl_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_wready = s_axi_control_wready;
end
always_comb begin // combinatorial s_axi_control_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bresp = 2'bxx;
	s_axi_control_bresp = _ctrl_bresp;
end
always_comb begin // combinatorial s_axi_control_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bvalid = 1'bx;
	s_axi_control_bvalid = _ctrl_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_bvalid = s_axi_control_bvalid;
end
always_comb begin // combinatorial s_axi_control_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_arready = 1'bx;
	s_axi_control_arready = _ctrl_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_arready = s_axi_control_arready;
end
always_comb begin // combinatorial s_axi_control_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	s_axi_control_rdata = _ctrl_rdata;
end
always_comb begin // combinatorial s_axi_control_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rresp = 2'bxx;
	s_axi_control_rresp = _ctrl_rresp;
end
always_comb begin // combinatorial s_axi_control_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rvalid = 1'bx;
	s_axi_control_rvalid = _ctrl_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_rvalid = s_axi_control_rvalid;
end
always_comb begin // combinatorial _ctrl_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awaddr = 12'dx;
	_ctrl_awaddr = s_axi_control_awaddr;
end
always_comb begin // combinatorial _ctrl_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awvalid = 1'bx;
	_ctrl_awvalid = s_axi_control_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_awvalid = _ctrl_awvalid;
end
always_comb begin // combinatorial _ctrl_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_ctrl_wdata = s_axi_control_wdata;
end
always_comb begin // combinatorial _ctrl_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wstrb = 4'bxxxx;
	_ctrl_wstrb = s_axi_control_wstrb;
end
always_comb begin // combinatorial _ctrl_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wvalid = 1'bx;
	_ctrl_wvalid = s_axi_control_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_wvalid = _ctrl_wvalid;
end
always_comb begin // combinatorial _ctrl_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_bready = 1'bx;
	_ctrl_bready = s_axi_control_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_bready = _ctrl_bready;
end
always_comb begin // combinatorial _ctrl_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_araddr = 12'dx;
	_ctrl_araddr = s_axi_control_araddr;
end
always_comb begin // combinatorial _ctrl_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_arvalid = 1'bx;
	_ctrl_arvalid = s_axi_control_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_arvalid = _ctrl_arvalid;
end
always_comb begin // combinatorial _ctrl_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_rready = 1'bx;
	_ctrl_rready = s_axi_control_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_rready = _ctrl_rready;
end
always_comb begin // combinatorial _reader_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_aresetn = 1'bx;
	_reader_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_aresetn = _reader_aresetn;
end
always_comb begin // combinatorial _writer_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_aresetn = 1'bx;
	_writer_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_aresetn = _writer_aresetn;
end
always_comb begin // combinatorial m_axi_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awvalid = 1'bx;
	m_axi_awvalid = _writer_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_awvalid = m_axi_awvalid;
end
always_comb begin // combinatorial m_axi_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awaddr = 64'dx;
	m_axi_awaddr = _writer_awaddr;
end
always_comb begin // combinatorial m_axi_awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awlen = 8'dx;
	m_axi_awlen = _writer_awlen;
end
always_comb begin // combinatorial m_axi_awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awburst = 2'bxx;
	m_axi_awburst = _writer_awburst;
end
always_comb begin // combinatorial m_axi_awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awcache = 4'bxxxx;
	m_axi_awcache = _writer_awcache;
end
always_comb begin // combinatorial m_axi_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wvalid = 1'bx;
	m_axi_wvalid = _writer_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wvalid = m_axi_wvalid;
end
always_comb begin // combinatorial m_axi_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wdata = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	m_axi_wdata = _writer_wdata;
end
always_comb begin // combinatorial m_axi_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wstrb = 8'bxxxxxxxx;
	m_axi_wstrb = _writer_wstrb;
end
always_comb begin // combinatorial m_axi_wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wlast = 1'bx;
	m_axi_wlast = _writer_wlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wlast = m_axi_wlast;
end
always_comb begin // combinatorial m_axi_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_bready = 1'bx;
	m_axi_bready = _writer_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_bready = m_axi_bready;
end
always_comb begin // combinatorial _writer_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_awready = 1'bx;
	_writer_awready = m_axi_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_awready = _writer_awready;
end
always_comb begin // combinatorial _writer_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_wready = 1'bx;
	_writer_wready = m_axi_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_wready = _writer_wready;
end
always_comb begin // combinatorial _writer_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bvalid = 1'bx;
	_writer_bvalid = m_axi_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_bvalid = _writer_bvalid;
end
always_comb begin // combinatorial _writer_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bresp = 2'bxx;
	_writer_bresp = m_axi_bresp;
end
always_comb begin // combinatorial m_axi_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arvalid = 1'bx;
	m_axi_arvalid = _reader_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arvalid = m_axi_arvalid;
end
always_comb begin // combinatorial m_axi_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_araddr = 64'dx;
	m_axi_araddr = _reader_araddr;
end
always_comb begin // combinatorial m_axi_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlen = 8'dx;
	m_axi_arlen = _reader_arlen;
end
always_comb begin // combinatorial m_axi_arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arsize = 3'dx;
	m_axi_arsize = _reader_arsize;
end
always_comb begin // combinatorial m_axi_arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arburst = 2'bxx;
	m_axi_arburst = _reader_arburst;
end
always_comb begin // combinatorial m_axi_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_rready = 1'bx;
	m_axi_rready = _reader_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_rready = m_axi_rready;
end
always_comb begin // combinatorial _reader_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_arready = 1'bx;
	_reader_arready = m_axi_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_arready = _reader_arready;
end
always_comb begin // combinatorial _reader_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rvalid = 1'bx;
	_reader_rvalid = m_axi_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rvalid = _reader_rvalid;
end
always_comb begin // combinatorial _reader_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rdata = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_reader_rdata = m_axi_rdata;
end
always_comb begin // combinatorial _reader_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rresp = 2'bxx;
	_reader_rresp = m_axi_rresp;
end
always_comb begin // combinatorial _reader_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rlast = 1'bx;
	_reader_rlast = m_axi_rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rlast = _reader_rlast;
end
always_comb begin // combinatorial addr_a_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	addr_a_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[_v0] = _46[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[32 + _v0] = _47[_v0];
end
end
always_comb begin // combinatorial start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	start_addr = 64'dx;
	start_addr = _BitsToUInt_value;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_BitsToUInt_bits = addr_a_bits;
end
always_comb begin // combinatorial num_to_transfer
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_to_transfer = 32'dx;
	num_to_transfer = _IntNarrow_out;
end
always_comb begin // combinatorial _BitsToUInt_2_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_2_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_BitsToUInt_2_bits = _49;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 32'dx;
	_IntNarrow_in = _BitsToUInt_2_value;
end
always_comb begin // combinatorial config_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	config_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	config_bits = _50;
end
always_comb begin // combinatorial m_axi_arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arprot = 3'bxxx;
	m_axi_arprot = _51;
end
always_comb begin // combinatorial m_axi_arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arcache = 4'bxxxx;
	m_axi_arcache = _52;
end
always_comb begin // combinatorial m_axi_arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arqos = 4'dx;
	m_axi_arqos = _BitsToUInt_3_value;
end
always_comb begin // combinatorial _BitsToUInt_3_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_3_bits = 4'bxxxx;
	_BitsToUInt_3_bits = _53;
end
always_comb begin // combinatorial m_axi_arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlock = 1'bx;
	m_axi_arlock = _54;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arlock = m_axi_arlock;
end
always_comb begin // combinatorial m_axi_arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arregion = 4'dx;
	m_axi_arregion = _BitsToUInt_4_value;
end
always_comb begin // combinatorial _BitsToUInt_4_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_4_bits = 4'bxxxx;
	_BitsToUInt_4_bits = _55;
end
always_comb begin // combinatorial _BitsToUInt_5_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_5_bits = 11'bxxxxxxxxxxx;
	_BitsToUInt_5_bits = _56;
end
always_comb begin // combinatorial _reader_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_max_in_flight = 11'dx;
	_reader_max_in_flight = _BitsToUInt_5_value;
end
always_ff @(posedge aclk) begin // state cycles_since_reset
	cycles_since_reset <= _60;
	if(_153) cycles_since_reset <= 1'd0;
end
always_comb begin // combinatorial cycles_since_reset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cycles_since_reset_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	cycles_since_reset_bits = __UIntToBits_bits_D3;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 64'dx;
	_UIntToBits_value = cycles_since_reset;
end
always_ff @(posedge aclk) begin // state cycles_since_reset_at_start
	if(__ctrl_start_D3) cycles_since_reset_at_start <= cycles_since_reset_bits;
end
always_ff @(posedge aclk) begin // state running
	if(_ctrl_start) running <= 1'b1;
	if(_reader_value_valid) if(last) running <= 1'b0;
	if(_153) running <= 1'b0;
end
always_ff @(posedge aclk) begin // state num_cycles_running
	if(_ctrl_start) num_cycles_running <= 1'd0;
	if(running) num_cycles_running <= _73;
	if(_153) num_cycles_running <= 1'd0;
end
always_ff @(posedge aclk) begin // state hash
	if(__ctrl_start_D2) hash <= _67;
	if(__reader_value_valid_D2) hash <= new_hash;
	if(__153_D2) hash <= _155;
end
always_comb begin // combinatorial _reader_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_request_new_burst = 1'bx;
	_reader_request_new_burst = 1'b0;
	if(_ctrl_start) _reader_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_request_new_burst = _reader_request_new_burst;
end
always_comb begin // combinatorial _reader_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_start_addr = 64'dx;
	if(_ctrl_start) _reader_start_addr = start_addr;
end
always_comb begin // combinatorial _reader_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_count = 32'dx;
	if(_ctrl_start) _reader_count = num_to_transfer;
end
always_comb begin // combinatorial _reader_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_is_ready_to_receive_lots_of_data = 1'bx;
	_reader_is_ready_to_receive_lots_of_data = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_is_ready_to_receive_lots_of_data = _reader_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
if(_reader_value_valid) value[_v0] = _reader_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_reader_value_valid) last = _reader_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_comb begin // combinatorial new_hash_contrib
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_hash_contrib = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(__reader_value_valid_D2) new_hash_contrib[0] = __75_D2;
	if(__reader_value_valid_D2) new_hash_contrib[1] = __77_D2;
	if(__reader_value_valid_D2) new_hash_contrib[2] = __79_D2;
	if(__reader_value_valid_D2) new_hash_contrib[3] = __81_D2;
	if(__reader_value_valid_D2) new_hash_contrib[4] = __83_D2;
	if(__reader_value_valid_D2) new_hash_contrib[5] = __85_D2;
	if(__reader_value_valid_D2) new_hash_contrib[6] = __87_D2;
	if(__reader_value_valid_D2) new_hash_contrib[7] = __89_D2;
	if(__reader_value_valid_D2) new_hash_contrib[8] = __91_D2;
	if(__reader_value_valid_D2) new_hash_contrib[9] = __93_D2;
	if(__reader_value_valid_D2) new_hash_contrib[10] = __95_D2;
	if(__reader_value_valid_D2) new_hash_contrib[11] = __97_D2;
	if(__reader_value_valid_D2) new_hash_contrib[12] = __99_D2;
	if(__reader_value_valid_D2) new_hash_contrib[13] = __101_D2;
	if(__reader_value_valid_D2) new_hash_contrib[14] = __103_D2;
	if(__reader_value_valid_D2) new_hash_contrib[15] = __105_D2;
	if(__reader_value_valid_D2) new_hash_contrib[16] = __107_D2;
	if(__reader_value_valid_D2) new_hash_contrib[17] = __109_D2;
	if(__reader_value_valid_D2) new_hash_contrib[18] = __111_D2;
	if(__reader_value_valid_D2) new_hash_contrib[19] = __113_D2;
	if(__reader_value_valid_D2) new_hash_contrib[20] = __115_D2;
	if(__reader_value_valid_D2) new_hash_contrib[21] = __117_D2;
	if(__reader_value_valid_D2) new_hash_contrib[22] = __119_D2;
	if(__reader_value_valid_D2) new_hash_contrib[23] = __121_D2;
	if(__reader_value_valid_D2) new_hash_contrib[24] = __123_D2;
	if(__reader_value_valid_D2) new_hash_contrib[25] = __125_D2;
	if(__reader_value_valid_D2) new_hash_contrib[26] = __127_D2;
	if(__reader_value_valid_D2) new_hash_contrib[27] = __129_D2;
	if(__reader_value_valid_D2) new_hash_contrib[28] = __131_D2;
	if(__reader_value_valid_D2) new_hash_contrib[29] = __133_D2;
	if(__reader_value_valid_D2) new_hash_contrib[30] = __135_D2;
	if(__reader_value_valid_D2) new_hash_contrib[31] = __137_D2;
end
always_comb begin // combinatorial new_hash
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_hash = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(__reader_value_valid_D2) new_hash = _140;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 32'dx;
	if(_reader_value_valid) if(last) _UIntToBits_2_value = num_cycles_running;
end
always_comb begin // combinatorial _ctrl_finish
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_finish = 1'bx;
	_ctrl_finish = 1'b0;
	if(__reader_value_valid_D3) if(_last_D3) _ctrl_finish = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_finish = _ctrl_finish;
end
always_comb begin // combinatorial _ctrl_output_regs
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_output_regs = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
if(__reader_value_valid_D3) if(_last_D3) _ctrl_output_regs[_v0] = _148[_v0];
end
end
endmodule

// axi_memory_writer_tie_off #(AXI_WIDTH: 64)
module axi_memory_writer_tie_off_AXI_WIDTH_64(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic awvalid,
	input wire awready,
	output /*mux_wire*/ logic[63:0] awaddr,
	output /*mux_wire*/ logic[7:0] awlen,
	output /*mux_wire*/ logic[2:0] awsize,
	output /*mux_wire*/ logic[1:0] awburst,
	output /*mux_wire*/ logic[2:0] awprot,
	output /*mux_wire*/ logic[3:0] awcache,
	output /*mux_wire*/ logic[3:0] awqos,
	output /*mux_wire*/ logic awlock,
	output /*mux_wire*/ logic[3:0] awregion,
	output /*mux_wire*/ logic wvalid,
	input wire wready,
	output /*mux_wire*/ logic[63:0] wdata,
	output /*mux_wire*/ logic[7:0] wstrb,
	output /*mux_wire*/ logic wlast,
	input wire bvalid,
	input wire[1:0] bresp,
	output /*mux_wire*/ logic bready
);

/*mux_wire*/ logic _aresetn;
localparam[1:0] _4 = 2'b00;
localparam[2:0] _5 = 3'b000;
localparam[3:0] _6 = 4'b0000;
/*mux_wire*/ logic _Repeat_v;
wire[63:0] _Repeat_result;
/*mux_wire*/ logic _Repeat_2_v;
wire[7:0] _Repeat_2_result;
/*mux_wire*/ logic _awready;
/*mux_wire*/ logic _wready;
/*mux_wire*/ logic _bvalid;
/*mux_wire*/ logic[1:0] _bresp;
Repeat_T_type_bool_SIZE_64 Repeat(
	.clk(aclk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
Repeat_T_type_bool_SIZE_8 Repeat_2(
	.clk(aclk),
	.v(_Repeat_2_v),
	.result(_Repeat_2_result)
);
always_comb begin // combinatorial _aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_aresetn = 1'bx;
	_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_aresetn = _aresetn;
end
always_comb begin // combinatorial awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awvalid = 1'bx;
	awvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awvalid = awvalid;
end
always_comb begin // combinatorial awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awaddr = 64'dx;
	awaddr = 1'd0;
end
always_comb begin // combinatorial awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlen = 8'dx;
	awlen = 1'd0;
end
always_comb begin // combinatorial awsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awsize = 3'dx;
	awsize = 2'd3;
end
always_comb begin // combinatorial awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awburst = 2'bxx;
	awburst = _4;
end
always_comb begin // combinatorial awprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awprot = 3'bxxx;
	awprot = _5;
end
always_comb begin // combinatorial awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awcache = 4'bxxxx;
	awcache = _6;
end
always_comb begin // combinatorial awqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awqos = 4'dx;
	awqos = 1'd0;
end
always_comb begin // combinatorial awlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlock = 1'bx;
	awlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awlock = awlock;
end
always_comb begin // combinatorial awregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awregion = 4'dx;
	awregion = 1'd0;
end
always_comb begin // combinatorial wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wvalid = 1'bx;
	wvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wvalid = wvalid;
end
always_comb begin // combinatorial wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wdata = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	wdata = _Repeat_result;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	_Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
always_comb begin // combinatorial wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wstrb = 8'bxxxxxxxx;
	wstrb = _Repeat_2_result;
end
always_comb begin // combinatorial _Repeat_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_2_v = 1'bx;
	_Repeat_2_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_2_v = _Repeat_2_v;
end
always_comb begin // combinatorial wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wlast = 1'bx;
	wlast = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wlast = wlast;
end
always_comb begin // combinatorial bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	bready = 1'bx;
	bready = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	bready = bready;
end
always_comb begin // combinatorial _awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_awready = 1'bx;
	_awready = awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_awready = _awready;
end
always_comb begin // combinatorial _wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_wready = 1'bx;
	_wready = wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_wready = _wready;
end
always_comb begin // combinatorial _bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_bvalid = 1'bx;
	_bvalid = bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_bvalid = _bvalid;
end
always_comb begin // combinatorial _bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_bresp = 2'bxx;
	_bresp = bresp;
end
endmodule

// Repeat #(T: type bool #(), SIZE: 8)
module Repeat_T_type_bool_SIZE_8(
	input clk,
	input wire v,
	output /*mux_wire*/ logic[7:0] result
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = 8'bxxxxxxxx;
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
	result[4] = v;
	result[5] = v;
	result[6] = v;
	result[7] = v;
end
endmodule

// Repeat #(T: type bool #(), SIZE: 64)
module Repeat_T_type_bool_SIZE_64(
	input clk,
	input wire v,
	output /*mux_wire*/ logic[63:0] result
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
	result[4] = v;
	result[5] = v;
	result[6] = v;
	result[7] = v;
	result[8] = v;
	result[9] = v;
	result[10] = v;
	result[11] = v;
	result[12] = v;
	result[13] = v;
	result[14] = v;
	result[15] = v;
	result[16] = v;
	result[17] = v;
	result[18] = v;
	result[19] = v;
	result[20] = v;
	result[21] = v;
	result[22] = v;
	result[23] = v;
	result[24] = v;
	result[25] = v;
	result[26] = v;
	result[27] = v;
	result[28] = v;
	result[29] = v;
	result[30] = v;
	result[31] = v;
	result[32] = v;
	result[33] = v;
	result[34] = v;
	result[35] = v;
	result[36] = v;
	result[37] = v;
	result[38] = v;
	result[39] = v;
	result[40] = v;
	result[41] = v;
	result[42] = v;
	result[43] = v;
	result[44] = v;
	result[45] = v;
	result[46] = v;
	result[47] = v;
	result[48] = v;
	result[49] = v;
	result[50] = v;
	result[51] = v;
	result[52] = v;
	result[53] = v;
	result[54] = v;
	result[55] = v;
	result[56] = v;
	result[57] = v;
	result[58] = v;
	result[59] = v;
	result[60] = v;
	result[61] = v;
	result[62] = v;
	result[63] = v;
end
endmodule

// axi_realigning_burst_reader #(T: type bool #()[32][2], AXI_WIDTH: 64, ADDR_ALIGN: 4, COUNT_TO: 4294967296, ATO: 18446744073709551616)
module axi_realigning_burst_reader_T_type_bool_32_2_AXI_WIDTH_64_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic arvalid,
	input wire arready,
	output /*mux_wire*/ logic[63:0] araddr,
	output /*mux_wire*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[63:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[31:0] count,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic value_valid,
	output /*mux_wire*/ logic[31:0] value[1:0],
	output /*mux_wire*/ logic last
);

/*mux_wire*/ logic _parent_aresetn;
wire _parent_arvalid;
wire[63:0] _parent_araddr;
wire[7:0] _parent_arlen;
wire[2:0] _parent_arsize;
wire[1:0] _parent_arburst;
wire[2:0] _parent_arprot;
wire[3:0] _parent_arcache;
wire[3:0] _parent_arqos;
wire _parent_arlock;
wire[3:0] _parent_arregion;
wire _parent_rready;
/*mux_wire*/ logic _parent_arready;
/*mux_wire*/ logic _parent_rvalid;
/*mux_wire*/ logic[63:0] _parent_rdata;
/*mux_wire*/ logic[1:0] _parent_rresp;
/*mux_wire*/ logic _parent_rlast;
/*mux_wire*/ logic[10:0] _parent_max_in_flight;
wire _parent_may_request_new_burst;
wire[32:0] _22;
assign _22 = count * 2'd2;
/*mux_wire*/ logic _parent_request_new_burst;
/*mux_wire*/ logic[63:0] _parent_start_addr;
/*mux_wire*/ logic[32:0] _parent_count;
/*mux_wire*/ logic _parent_is_ready_to_receive_lots_of_data;
/*state*/ logic[31:0] stored_elements[0:0];
/*state*/ logic[0:0] cur_element_store_align;
wire _parent_element_packet_valid;
wire[31:0] _parent_elements[1:0];
wire[0:0] _parent_chunk_offset;
wire[1:0] _parent_chunk_length;
wire _parent_last;
/*mux_wire*/ logic[31:0] elements[1:0];
/*mux_wire*/ logic[0:0] chunk_offset;
/*mux_wire*/ logic[1:0] chunk_length;
/*mux_wire*/ logic last_2;
/*mux_wire*/ logic[31:0] elements_extended[1:0];
/*mux_wire*/ logic[31:0] rotated_elements[1:0];
wire signed[1:0] _31;
assign _31 = cur_element_store_align - chunk_offset;
wire[0:0] _32;
assign _32 = _31; // == mod 2 (target is 1 bits wide)
/*mux_wire*/ logic[31:0] _RotateRight_data[1:0];
/*mux_wire*/ logic[0:0] _RotateRight_offset;
wire[31:0] _RotateRight_rotated_data[1:0];
/*mux_wire*/ logic[1:0] rotated_strobe;
/*mux_wire*/ logic[0:0] _MakeStrobe_chunk_offset;
/*mux_wire*/ logic[1:0] _MakeStrobe_chunk_length;
wire[1:0] _MakeStrobe_strobe;
/*mux_wire*/ logic[1:0] end_of_element;
wire[1:0] _37;
assign _37 = cur_element_store_align + chunk_length;
wire _39;
assign _39 = end_of_element >= 2'd2;
/*mux_wire*/ logic[63:0] resulting_value_bits;
wire _41;
assign _41 = cur_element_store_align > 1'd0;
wire[31:0] _42 = stored_elements[0];
wire[31:0] _43 = rotated_elements[0];
wire[31:0] _44 = rotated_elements[1];
/*mux_wire*/ logic[63:0] _FromBits_bits;
wire[31:0] _FromBits_value[1:0];
wire[0:0] _49;
assign _49 = end_of_element; // == mod 2 (target is 1 bits wide)
wire _50 = rotated_strobe[0];
wire[31:0] _51 = rotated_elements[0];
wire _53;
assign _53 = !aresetn;
axi_array_burst_reader_AXI_WIDTH_64_ADDR_ALIGN_4_COUNT_TO_8589934592_ATO_18446744073709551616 parent(
	.aclk(aclk),
	.aresetn(_parent_aresetn),
	.arvalid(_parent_arvalid),
	.arready(_parent_arready),
	.araddr(_parent_araddr),
	.arlen(_parent_arlen),
	.arsize(_parent_arsize),
	.arburst(_parent_arburst),
	.arprot(_parent_arprot),
	.arcache(_parent_arcache),
	.arqos(_parent_arqos),
	.arlock(_parent_arlock),
	.arregion(_parent_arregion),
	.rvalid(_parent_rvalid),
	.rready(_parent_rready),
	.rdata(_parent_rdata),
	.rresp(_parent_rresp),
	.rlast(_parent_rlast),
	.is_ready_to_receive_lots_of_data(_parent_is_ready_to_receive_lots_of_data),
	.element_packet_valid(_parent_element_packet_valid),
	.elements(_parent_elements),
	.chunk_offset(_parent_chunk_offset),
	.chunk_length(_parent_chunk_length),
	.last(_parent_last),
	.max_in_flight(_parent_max_in_flight),
	.may_request_new_burst(_parent_may_request_new_burst),
	.request_new_burst(_parent_request_new_burst),
	.start_addr(_parent_start_addr),
	.count(_parent_count)
);
RotateRight_T_type_bool_32_ARRAY_LEN_2 RotateRight(
	.clk(aclk),
	.data(_RotateRight_data),
	.offset(_RotateRight_offset),
	.rotated_data(_RotateRight_rotated_data)
);
MakeStrobe_STROBE_WIDTH_2 MakeStrobe(
	.clk(aclk),
	.chunk_offset(_MakeStrobe_chunk_offset),
	.chunk_length(_MakeStrobe_chunk_length),
	.strobe(_MakeStrobe_strobe)
);
FromBits_T_type_bool_32_2 FromBits(
	.clk(aclk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial _parent_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_aresetn = 1'bx;
	_parent_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_aresetn = _parent_aresetn;
end
always_comb begin // combinatorial arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arvalid = 1'bx;
	arvalid = _parent_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arvalid = arvalid;
end
always_comb begin // combinatorial araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	araddr = 64'dx;
	araddr = _parent_araddr;
end
always_comb begin // combinatorial arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlen = 8'dx;
	arlen = _parent_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = _parent_arsize;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _parent_arburst;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _parent_arprot;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _parent_arcache;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = _parent_arqos;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = _parent_arlock;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = _parent_arregion;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = _parent_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _parent_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_arready = 1'bx;
	_parent_arready = arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_arready = _parent_arready;
end
always_comb begin // combinatorial _parent_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rvalid = 1'bx;
	_parent_rvalid = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rvalid = _parent_rvalid;
end
always_comb begin // combinatorial _parent_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rdata = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_parent_rdata = rdata;
end
always_comb begin // combinatorial _parent_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rresp = 2'bxx;
	_parent_rresp = rresp;
end
always_comb begin // combinatorial _parent_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rlast = 1'bx;
	_parent_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rlast = _parent_rlast;
end
always_comb begin // combinatorial _parent_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_max_in_flight = 11'dx;
	_parent_max_in_flight = max_in_flight;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _parent_may_request_new_burst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial _parent_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_request_new_burst = 1'bx;
	_parent_request_new_burst = 1'b0;
	if(request_new_burst) _parent_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_request_new_burst = _parent_request_new_burst;
end
always_comb begin // combinatorial _parent_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_start_addr = 64'dx;
	if(request_new_burst) _parent_start_addr = start_addr;
end
always_comb begin // combinatorial _parent_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_count = 33'dx;
	if(request_new_burst) _parent_count = _22;
end
always_comb begin // combinatorial _parent_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_is_ready_to_receive_lots_of_data = 1'bx;
	_parent_is_ready_to_receive_lots_of_data = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_is_ready_to_receive_lots_of_data = _parent_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value_valid = 1'bx;
	value_valid = 1'b0;
	if(_parent_element_packet_valid) if(_39) value_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	value_valid = value_valid;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) value[_v0] = _FromBits_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_parent_element_packet_valid) if(_39) last = last_2;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state stored_elements
	if(_parent_element_packet_valid) if(_50) stored_elements[0] <= _51;
end
always_ff @(posedge aclk) begin // state cur_element_store_align
	if(_parent_element_packet_valid) cur_element_store_align <= _49;
	if(_53) cur_element_store_align <= 1'd0;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements[_v0] = _parent_elements[_v0];
end
end
always_comb begin // combinatorial chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_offset = 1'dx;
	if(_parent_element_packet_valid) chunk_offset = _parent_chunk_offset;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunk_offset = chunk_offset;
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 2'dx;
	if(_parent_element_packet_valid) chunk_length = _parent_chunk_length;
end
always_comb begin // combinatorial last_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last_2 = 1'bx;
	if(_parent_element_packet_valid) last_2 = _parent_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last_2 = last_2;
end
always_comb begin // combinatorial elements_extended
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_extended = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements_extended[_v0] = elements[_v0];
end
end
always_comb begin // combinatorial rotated_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) rotated_elements[_v0] = _RotateRight_rotated_data[_v0];
end
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) _RotateRight_data[_v0] = elements_extended[_v0];
end
end
always_comb begin // combinatorial _RotateRight_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_offset = 1'dx;
	if(_parent_element_packet_valid) _RotateRight_offset = _32;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_RotateRight_offset = _RotateRight_offset;
end
always_comb begin // combinatorial rotated_strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_strobe = 2'bxx;
	if(_parent_element_packet_valid) rotated_strobe = _MakeStrobe_strobe;
end
always_comb begin // combinatorial _MakeStrobe_chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_offset = 1'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_offset = cur_element_store_align;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_MakeStrobe_chunk_offset = _MakeStrobe_chunk_offset;
end
always_comb begin // combinatorial _MakeStrobe_chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_length = 2'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_length = chunk_length;
end
always_comb begin // combinatorial end_of_element
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	end_of_element = 2'dx;
	if(_parent_element_packet_valid) end_of_element = _37;
end
always_comb begin // combinatorial resulting_value_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	resulting_value_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_41) resulting_value_bits[_v0] = _42[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_41) resulting_value_bits[_v0] = _43[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) resulting_value_bits[32 + _v0] = _44[_v0];
end
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_parent_element_packet_valid) if(_39) _FromBits_bits = resulting_value_bits;
end
endmodule

// FromBits #(T: type bool #()[32][2])
module FromBits_T_type_bool_32_2(
	input clk,
	input wire[63:0] bits,
	output /*mux_wire*/ logic[31:0] value[1:0]
);

genvar _g0;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign value[_g0] = bits[(_g0) * 32 +: 32];
end
endgenerate
endmodule

// MakeStrobe #(STROBE_WIDTH: 2)
module MakeStrobe_STROBE_WIDTH_2(
	input clk,
	input wire[0:0] chunk_offset,
	input wire[1:0] chunk_length,
	output /*mux_wire*/ logic[1:0] strobe
);

/*mux_wire*/ logic[1:0] chunk_bits;
wire _2;
assign _2 = chunk_length > 1'd0;
wire _4;
assign _4 = chunk_length > 1'd1;
/*mux_wire*/ logic[1:0] _RotateRight_data;
/*mux_wire*/ logic[0:0] _RotateRight_offset;
wire[1:0] _RotateRight_rotated_data;
RotateRight_T_type_bool_ARRAY_LEN_2 RotateRight(
	.clk(clk),
	.data(_RotateRight_data),
	.offset(_RotateRight_offset),
	.rotated_data(_RotateRight_rotated_data)
);
always_comb begin // combinatorial strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	strobe = 2'bxx;
	strobe = _RotateRight_rotated_data;
end
always_comb begin // combinatorial chunk_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_bits = 2'bxx;
	if(_2) chunk_bits[0] = 1'b1;
	if(!_2) chunk_bits[0] = 1'b0;
	if(_4) chunk_bits[1] = 1'b1;
	if(!_4) chunk_bits[1] = 1'b0;
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = 2'bxx;
	_RotateRight_data = chunk_bits;
end
always_comb begin // combinatorial _RotateRight_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_offset = 1'dx;
	_RotateRight_offset = chunk_offset;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_RotateRight_offset = _RotateRight_offset;
end
endmodule

// RotateRight #(T: type bool #(), ARRAY_LEN: 2)
module RotateRight_T_type_bool_ARRAY_LEN_2(
	input clk,
	input wire[1:0] data,
	input wire[0:0] offset,
	output /*mux_wire*/ logic[1:0] rotated_data
);

/*mux_wire*/ logic[0:0] offset_bits;
/*mux_wire*/ logic[0:0] _UIntToBits_value;
wire[0:0] _UIntToBits_bits;
/*mux_wire*/ logic[1:0] rotate_stages[1:0];
/*mux_wire*/ logic[1:0] from;
wire[1:0] _3 = rotate_stages[0];
wire _4 = offset_bits[0];
wire _5 = from[1];
wire _6 = from[0];
wire _7 = offset_bits[0];
wire _8 = from[0];
wire _9 = from[1];
wire[1:0] _10 = rotate_stages[1];
UIntToBits_NUM_BITS_1 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = 2'bxx;
	rotated_data = _10;
end
always_comb begin // combinatorial offset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	offset_bits = 1'bx;
	offset_bits = _UIntToBits_bits;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	offset_bits = offset_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 1'dx;
	_UIntToBits_value = offset;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_UIntToBits_value = _UIntToBits_value;
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{2'bxx, 2'bxx};
	rotate_stages[0] = data;
	if(_4) rotate_stages[1][0] = _5;
	if(!_4) rotate_stages[1][0] = _6;
	if(_7) rotate_stages[1][1] = _8;
	if(!_7) rotate_stages[1][1] = _9;
end
always_comb begin // combinatorial from
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from = 2'bxx;
	from = _3;
end
endmodule

// RotateRight #(T: type bool #()[32], ARRAY_LEN: 2)
module RotateRight_T_type_bool_32_ARRAY_LEN_2(
	input clk,
	input wire[31:0] data[1:0],
	input wire[0:0] offset,
	output /*mux_wire*/ logic[31:0] rotated_data[1:0]
);

genvar _g0;
/*mux_wire*/ logic[0:0] offset_bits;
/*mux_wire*/ logic[0:0] _UIntToBits_value;
wire[0:0] _UIntToBits_bits;
/*mux_wire*/ logic[31:0] rotate_stages[1:0][1:0];
/*mux_wire*/ logic[31:0] from[1:0];
wire[31:0] _3[1:0];
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _3[_g0] = rotate_stages[0][_g0];
end
endgenerate
wire _4 = offset_bits[0];
wire[31:0] _5 = from[1];
wire[31:0] _6 = from[0];
wire _7 = offset_bits[0];
wire[31:0] _8 = from[0];
wire[31:0] _9 = from[1];
wire[31:0] _10[1:0];
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _10[_g0] = rotate_stages[1][_g0];
end
endgenerate
UIntToBits_NUM_BITS_1 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
rotated_data[_v0] = _10[_v0];
end
end
always_comb begin // combinatorial offset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	offset_bits = 1'bx;
	offset_bits = _UIntToBits_bits;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	offset_bits = offset_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 1'dx;
	_UIntToBits_value = offset;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_UIntToBits_value = _UIntToBits_value;
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{'{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}};
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
rotate_stages[0][_v0] = data[_v0];
end
	if(_4) rotate_stages[1][0] = _5;
	if(!_4) rotate_stages[1][0] = _6;
	if(_7) rotate_stages[1][1] = _8;
	if(!_7) rotate_stages[1][1] = _9;
end
always_comb begin // combinatorial from
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
from[_v0] = _3[_v0];
end
end
endmodule

// axi_array_burst_reader #(AXI_WIDTH: 64, ADDR_ALIGN: 4, COUNT_TO: 8589934592, ATO: 18446744073709551616)
module axi_array_burst_reader_AXI_WIDTH_64_ADDR_ALIGN_4_COUNT_TO_8589934592_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*state*/ logic arvalid,
	input wire arready,
	output /*state*/ logic[63:0] araddr,
	output /*state*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[63:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic element_packet_valid,
	output /*mux_wire*/ logic[31:0] elements[1:0],
	output /*mux_wire*/ logic[0:0] chunk_offset,
	output /*mux_wire*/ logic[1:0] chunk_length,
	output /*mux_wire*/ logic last,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[32:0] count
);

/*latency*/ logic _arvalid_D1; always_ff @(posedge aclk) begin _arvalid_D1 <= arvalid; end
/*latency*/ logic _request_new_burst_D1; always_ff @(posedge aclk) begin _request_new_burst_D1 <= request_new_burst; end
genvar _g0;
localparam[1:0] _1 = 2'b01;
localparam[2:0] _2 = 3'b000;
localparam[3:0] _3 = 4'b0010;
/*mux_wire*/ logic[1:0] _rresp;
/*mux_wire*/ logic _rlast;
/*state*/ logic[11:0] num_in_flight;
/*state*/ logic last_burst_in_flight;
/*mux_wire*/ logic[63:0] next_araddr;
/*latency*/ logic[63:0] _next_araddr_D0; always_ff @(posedge aclk) begin _next_araddr_D0 <= next_araddr; end
wire[60:0] _cur_start_chunk_addr_old;
/*mux_wire*/ logic[60:0] _BitwiseIntConcat_upper;
/*mux_wire*/ logic[2:0] _BitwiseIntConcat_lower;
wire[63:0] _BitwiseIntConcat_v;
/*mux_wire*/ logic[7:0] next_arlen;
/*mux_wire*/ logic next_last_burst_in_flight;
/*latency*/ logic _next_last_burst_in_flight_D0; always_ff @(posedge aclk) begin _next_last_burst_in_flight_D0 <= next_last_burst_in_flight; end
/*mux_wire*/ logic[52:0] cur_burst_addr;
/*mux_wire*/ logic[7:0] cur_align;
/*mux_wire*/ logic[60:0] _BitwiseIntSplit_v;
wire[52:0] _BitwiseIntSplit_upper;
wire[7:0] _BitwiseIntSplit_lower;
/*mux_wire*/ logic chunks_are_left;
/*latency*/ logic _chunks_are_left_D0; always_ff @(posedge aclk) begin _chunks_are_left_D0 <= chunks_are_left; end
wire[32:0] _num_chunks_left_old;
/*latency*/ logic[32:0] __num_chunks_left_old_N1; always_ff @(posedge aclk) begin __num_chunks_left_old_N1 <= _num_chunks_left_old; end
/*latency*/ logic[32:0] __num_chunks_left_old_D0; always_ff @(posedge aclk) begin __num_chunks_left_old_D0 <= __num_chunks_left_old_N1; end
wire _14;
assign _14 = _num_chunks_left_old > 1'd0;
/*latency*/ logic __14_N1; always_ff @(posedge aclk) begin __14_N1 <= _14; end
/*mux_wire*/ logic[7:0] max_chunks_in_this_burst;
/*latency*/ logic[7:0] _max_chunks_in_this_burst_D0; always_ff @(posedge aclk) begin _max_chunks_in_this_burst_D0 <= max_chunks_in_this_burst; end
wire[7:0] _18;
assign _18 = 8'd255 - cur_align;
wire[8:0] _22;
assign _22 = max_chunks_in_this_burst + 1'd1;
wire _23;
assign _23 = __num_chunks_left_old_N1 <= _22;
/*latency*/ logic __23_D0; always_ff @(posedge aclk) begin __23_D0 <= _23; end
/*mux_wire*/ logic[32:0] _IntNarrow_in;
wire[8:0] _IntNarrow_out;
wire[7:0] _26;
assign _26 = _IntNarrow_out - 1'd1;
/*latency*/ logic[7:0] __26_D0; always_ff @(posedge aclk) begin __26_D0 <= _26; end
/*mux_wire*/ logic may_next_arvalid;
/*latency*/ logic _may_next_arvalid_D1; always_ff @(posedge aclk) begin _may_next_arvalid_D1 <= may_next_arvalid; end
wire _num_chunks_left_may_update;
wire _30;
assign _30 = _chunks_are_left_D0 & _num_chunks_left_may_update;
wire _cur_start_chunk_addr_may_update;
wire _32;
assign _32 = _30 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
wire _34;
assign _34 = _32 & _LatencyOffset_out;
wire signed[11:0] _37;
assign _37 = max_in_flight - 9'd256;
wire _38;
assign _38 = $signed({1'b0, num_in_flight}) <= _37;
wire _39;
assign _39 = _34 & _38;
/*mux_wire*/ logic[53:0] next_burst_addr;
wire[53:0] _45;
assign _45 = cur_burst_addr + 1'd1;
/*latency*/ logic[53:0] __45_D0; always_ff @(posedge aclk) begin __45_D0 <= _45; end
/*latency*/ logic[53:0] __45_D1; always_ff @(posedge aclk) begin __45_D1 <= __45_D0; end
/*mux_wire*/ logic[53:0] _BitwiseIntConcat_2_upper;
/*mux_wire*/ logic[7:0] _BitwiseIntConcat_2_lower;
wire[61:0] _BitwiseIntConcat_2_v;
/*mux_wire*/ logic[61:0] _IntNarrow_2_in;
wire[60:0] _IntNarrow_2_out;
/*mux_wire*/ logic _cur_start_chunk_addr_update;
/*mux_wire*/ logic[60:0] _cur_start_chunk_addr_new;
/*mux_wire*/ logic[32:0] next_num_chunks_left;
wire[8:0] _53;
assign _53 = next_arlen + 1'd1;
wire signed[33:0] _54;
assign _54 = __num_chunks_left_old_D0 - _53;
/*mux_wire*/ logic signed[33:0] _IntNarrow_3_in;
wire[32:0] _IntNarrow_3_out;
/*mux_wire*/ logic _num_chunks_left_update;
/*mux_wire*/ logic[32:0] _num_chunks_left_new;
/*mux_wire*/ logic _BoolToInt_i;
wire[0:0] _BoolToInt_o;
wire signed[12:0] _64;
assign _64 = num_in_flight - _BoolToInt_o;
wire _66;
assign _66 = !arvalid;
wire _68;
assign _68 = _66 & may_next_arvalid;
wire[8:0] _71;
assign _71 = next_arlen + 1'd1;
/*mux_wire*/ logic _Ternary_cond;
/*mux_wire*/ logic[8:0] _Ternary_a;
/*mux_wire*/ logic[8:0] _Ternary_b;
wire[8:0] _Ternary_o;
wire signed[12:0] _73;
assign _73 = _64 + $signed({1'b0, _Ternary_o});
/*mux_wire*/ logic signed[12:0] _IntNarrow_4_in;
wire[11:0] _IntNarrow_4_out;
/*state*/ logic[1:0] final_chunk_align;
/*state*/ logic[0:0] cur_chunk_align;
/*mux_wire*/ logic[31:0] elements_2[1:0];
wire[31:0] _75;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _75[_g0] = rdata[_g0];
end
endgenerate
wire[31:0] _76;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _76[_g0] = rdata[32 + _g0];
end
endgenerate
/*mux_wire*/ logic[1:0] num_chunk_elements;
/*mux_wire*/ logic is_last;
wire _79;
assign _79 = num_in_flight == 1'd1;
wire _81;
assign _81 = _79 & last_burst_in_flight;
wire signed[2:0] _85;
assign _85 = final_chunk_align - cur_chunk_align;
/*mux_wire*/ logic signed[2:0] _IntNarrow_5_in;
wire[1:0] _IntNarrow_5_out;
wire[1:0] _87;
assign _87 = 2'd2 - cur_chunk_align;
wire _95;
assign _95 = !chunks_are_left;
/*latency*/ logic __95_D0; always_ff @(posedge aclk) begin __95_D0 <= _95; end
wire _97;
assign _97 = __95_D0 & _num_chunks_left_may_update;
wire _99;
assign _99 = _97 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic[60:0] chunk_addr;
/*latency*/ logic[60:0] _chunk_addr_D1; always_ff @(posedge aclk) begin _chunk_addr_D1 <= chunk_addr; end
/*mux_wire*/ logic[0:0] element_in_chunk_align;
wire[61:0] _101;
assign _101 = start_addr / 3'd4;
/*mux_wire*/ logic[61:0] _BitwiseIntSplit_2_v;
wire[60:0] _BitwiseIntSplit_2_upper;
wire[0:0] _BitwiseIntSplit_2_lower;
/*mux_wire*/ logic[32:0] chunk_count_bits;
/*mux_wire*/ logic[0:0] final_alignment;
wire[33:0] _104;
assign _104 = count + element_in_chunk_align;
/*mux_wire*/ logic[33:0] _BitwiseIntSplit_3_v;
wire[32:0] _BitwiseIntSplit_3_upper;
wire[0:0] _BitwiseIntSplit_3_lower;
/*mux_wire*/ logic[32:0] num_chunks;
/*mux_wire*/ logic is_no_chunks;
wire _107;
assign _107 = chunk_count_bits == 1'd0;
wire _113;
assign _113 = final_alignment != 1'd0;
/*mux_wire*/ logic _BoolToInt_2_i;
wire[0:0] _BoolToInt_2_o;
wire[32:0] _114;
assign _114 = chunk_count_bits + _BoolToInt_2_o;
wire _120;
assign _120 = !is_no_chunks;
wire _123;
assign _123 = final_alignment == 1'd0;
wire _124;
assign _124 = _120 & _123;
/*mux_wire*/ logic _BoolToInt_3_i;
wire[0:0] _BoolToInt_3_o;
/*mux_wire*/ logic[0:0] _BitwiseIntConcat_3_upper;
/*mux_wire*/ logic[0:0] _BitwiseIntConcat_3_lower;
wire[1:0] _BitwiseIntConcat_3_v;
wire _128;
assign _128 = !aresetn;
/*mux_wire*/ logic _cur_start_chunk_addr_rst;
wire _130;
assign _130 = !aresetn;
/*mux_wire*/ logic _num_chunks_left_rst;
wire _132;
assign _132 = !aresetn;
SlowState_T_type_int_FROM_0_TO_2305843009213693952_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1 cur_start_chunk_addr(
	.clk(aclk),
	.rst(_cur_start_chunk_addr_rst),
	.old(_cur_start_chunk_addr_old),
	.may_update(_cur_start_chunk_addr_may_update),
	.update(_cur_start_chunk_addr_update),
	.new_1(_cur_start_chunk_addr_new)
);
SlowState_T_type_int_FROM_0_TO_4294967299_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0 num_chunks_left(
	.clk(aclk),
	.rst(_num_chunks_left_rst),
	.old(_num_chunks_left_old),
	.may_update(_num_chunks_left_may_update),
	.update(_num_chunks_left_update),
	.new_1(_num_chunks_left_new)
);
BitwiseIntConcat_UPPER_TO_2305843009213693952_LOWER_BITS_3 BitwiseIntConcat(
	.clk(aclk),
	.upper(_BitwiseIntConcat_upper),
	.lower(_BitwiseIntConcat_lower),
	.v(_BitwiseIntConcat_v)
);
BitwiseIntSplit_TO_2305843009213693952_LOWER_BITS_8 BitwiseIntSplit(
	.clk(aclk),
	.v(_BitwiseIntSplit_v),
	.upper(_BitwiseIntSplit_upper),
	.lower(_BitwiseIntSplit_lower)
);
IntNarrow_FROM_I_0_TO_I_4294967299_FROM_1_TO_257 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
LatencyOffset_T_type_bool_OFFSET_384 LatencyOffset(
	.clk(aclk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
BitwiseIntConcat_UPPER_TO_9007199254740993_LOWER_BITS_8 BitwiseIntConcat_2(
	.clk(aclk),
	.upper(_BitwiseIntConcat_2_upper),
	.lower(_BitwiseIntConcat_2_lower),
	.v(_BitwiseIntConcat_2_v)
);
IntNarrow_FROM_I_0_TO_I_2305843009213694208_FROM_0_TO_2305843009213693952 IntNarrow_2(
	.clk(aclk),
	.in(_IntNarrow_2_in),
	.out(_IntNarrow_2_out)
);
IntNarrow_FROM_I_256_TO_I_4294967298_FROM_0_TO_4294967299 IntNarrow_3(
	.clk(aclk),
	.in(_IntNarrow_3_in),
	.out(_IntNarrow_3_out)
);
BoolToInt BoolToInt(
	.clk(aclk),
	.i(_BoolToInt_i),
	.o(_BoolToInt_o)
);
Ternary_T_type_int_FROM_0_TO_257 Ternary(
	.clk(aclk),
	.cond(_Ternary_cond),
	.a(_Ternary_a),
	.b(_Ternary_b),
	.o(_Ternary_o)
);
IntNarrow_FROM_I_1_TO_I_3640_FROM_0_TO_3384 IntNarrow_4(
	.clk(aclk),
	.in(_IntNarrow_4_in),
	.out(_IntNarrow_4_out)
);
IntNarrow_FROM_I_1_TO_I_4_FROM_0_TO_3 IntNarrow_5(
	.clk(aclk),
	.in(_IntNarrow_5_in),
	.out(_IntNarrow_5_out)
);
BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_1 BitwiseIntSplit_2(
	.clk(aclk),
	.v(_BitwiseIntSplit_2_v),
	.upper(_BitwiseIntSplit_2_upper),
	.lower(_BitwiseIntSplit_2_lower)
);
BitwiseIntSplit_TO_8589934593_LOWER_BITS_1 BitwiseIntSplit_3(
	.clk(aclk),
	.v(_BitwiseIntSplit_3_v),
	.upper(_BitwiseIntSplit_3_upper),
	.lower(_BitwiseIntSplit_3_lower)
);
BoolToInt BoolToInt_2(
	.clk(aclk),
	.i(_BoolToInt_2_i),
	.o(_BoolToInt_2_o)
);
BoolToInt BoolToInt_3(
	.clk(aclk),
	.i(_BoolToInt_3_i),
	.o(_BoolToInt_3_o)
);
BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_1 BitwiseIntConcat_3(
	.clk(aclk),
	.upper(_BitwiseIntConcat_3_upper),
	.lower(_BitwiseIntConcat_3_lower),
	.v(_BitwiseIntConcat_3_v)
);
always_ff @(posedge aclk) begin // state arvalid
	if(arvalid) if(arready) arvalid <= 1'b0;
	if(!arvalid) if(may_next_arvalid) arvalid <= 1'b1;
	if(_132) arvalid <= 1'b0;
end
always_ff @(posedge aclk) begin // state araddr
	if(!arvalid) if(may_next_arvalid) araddr <= _next_araddr_D0;
end
always_ff @(posedge aclk) begin // state arlen
	if(!arvalid) if(may_next_arvalid) arlen <= next_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = 2'd3;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _1;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _2;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _3;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = 1'd0;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = 1'd0;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rresp = 2'bxx;
	_rresp = rresp;
end
always_comb begin // combinatorial _rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rlast = 1'bx;
	_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_rlast = _rlast;
end
always_comb begin // combinatorial element_packet_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_packet_valid = 1'bx;
	element_packet_valid = 1'b0;
	if(rvalid) element_packet_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	element_packet_valid = element_packet_valid;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
if(rvalid) elements[_v0] = elements_2[_v0];
end
end
always_comb begin // combinatorial chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_offset = 1'dx;
	if(rvalid) chunk_offset = cur_chunk_align;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunk_offset = chunk_offset;
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 2'dx;
	if(rvalid) chunk_length = num_chunk_elements;
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(rvalid) last = is_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state num_in_flight
	num_in_flight <= _IntNarrow_4_out;
	if(_132) num_in_flight <= 1'd0;
end
always_ff @(posedge aclk) begin // state last_burst_in_flight
	if(!arvalid) if(may_next_arvalid) last_burst_in_flight <= _next_last_burst_in_flight_D0;
end
always_comb begin // combinatorial next_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_araddr = 64'dx;
	next_araddr = _BitwiseIntConcat_v;
end
always_comb begin // combinatorial _BitwiseIntConcat_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_upper = 61'dx;
	_BitwiseIntConcat_upper = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial _BitwiseIntConcat_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_lower = 3'dx;
	_BitwiseIntConcat_lower = 1'd0;
end
always_comb begin // combinatorial next_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_arlen = 8'dx;
	if(_chunks_are_left_D0) if(__23_D0) next_arlen = __26_D0;
	if(_chunks_are_left_D0) if(!__23_D0) next_arlen = _max_chunks_in_this_burst_D0;
end
always_comb begin // combinatorial next_last_burst_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_last_burst_in_flight = 1'bx;
	next_last_burst_in_flight = 1'b0;
	if(chunks_are_left) if(_23) next_last_burst_in_flight = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	next_last_burst_in_flight = next_last_burst_in_flight;
end
always_comb begin // combinatorial cur_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_burst_addr = 53'dx;
	cur_burst_addr = _BitwiseIntSplit_upper;
end
always_comb begin // combinatorial cur_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_align = 8'dx;
	cur_align = _BitwiseIntSplit_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_v = 61'dx;
	_BitwiseIntSplit_v = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial chunks_are_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunks_are_left = 1'bx;
	chunks_are_left = __14_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunks_are_left = chunks_are_left;
end
always_comb begin // combinatorial max_chunks_in_this_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	max_chunks_in_this_burst = 8'dx;
	if(chunks_are_left) max_chunks_in_this_burst = _18;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 33'dx;
	if(chunks_are_left) if(_23) _IntNarrow_in = __num_chunks_left_old_N1;
end
always_comb begin // combinatorial may_next_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_next_arvalid = 1'bx;
	may_next_arvalid = _39;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_next_arvalid = may_next_arvalid;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial next_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_burst_addr = 54'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) next_burst_addr = __45_D1;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_upper = 54'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_upper = next_burst_addr;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_lower = 8'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_lower = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_2_in = 62'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _IntNarrow_2_in = _BitwiseIntConcat_2_v;
end
always_comb begin // combinatorial _cur_start_chunk_addr_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_update = 1'bx;
	_cur_start_chunk_addr_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _cur_start_chunk_addr_update = 1'b1;
	if(request_new_burst) _cur_start_chunk_addr_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_update = _cur_start_chunk_addr_update;
end
always_comb begin // combinatorial _cur_start_chunk_addr_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_new = 61'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _cur_start_chunk_addr_new = _IntNarrow_2_out;
	if(_request_new_burst_D1) _cur_start_chunk_addr_new = _chunk_addr_D1;
end
always_comb begin // combinatorial next_num_chunks_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_num_chunks_left = 33'dx;
	if(!arvalid) if(may_next_arvalid) next_num_chunks_left = _IntNarrow_3_out;
end
always_comb begin // combinatorial _IntNarrow_3_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_3_in = 34'sdx;
	if(!arvalid) if(may_next_arvalid) _IntNarrow_3_in = _54;
end
always_comb begin // combinatorial _num_chunks_left_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_update = 1'bx;
	_num_chunks_left_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_update = 1'b1;
	if(request_new_burst) _num_chunks_left_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_update = _num_chunks_left_update;
end
always_comb begin // combinatorial _num_chunks_left_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_new = 33'dx;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_new = next_num_chunks_left;
	if(request_new_burst) _num_chunks_left_new = num_chunks;
end
always_comb begin // combinatorial _BoolToInt_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_i = 1'bx;
	_BoolToInt_i = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_i = _BoolToInt_i;
end
always_comb begin // combinatorial _Ternary_cond
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_cond = 1'bx;
	_Ternary_cond = _68;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Ternary_cond = _Ternary_cond;
end
always_comb begin // combinatorial _Ternary_a
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_a = 9'dx;
	_Ternary_a = _71;
end
always_comb begin // combinatorial _Ternary_b
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_b = 9'dx;
	_Ternary_b = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_4_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_4_in = 13'sdx;
	_IntNarrow_4_in = _73;
end
always_ff @(posedge aclk) begin // state final_chunk_align
	if(request_new_burst) final_chunk_align <= _BitwiseIntConcat_3_v;
end
always_ff @(posedge aclk) begin // state cur_chunk_align
	if(rvalid) cur_chunk_align <= 1'd0;
	if(request_new_burst) cur_chunk_align <= element_in_chunk_align;
end
always_comb begin // combinatorial elements_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_2 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	if(rvalid) elements_2[0] = _75;
	if(rvalid) elements_2[1] = _76;
end
always_comb begin // combinatorial num_chunk_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunk_elements = 2'dx;
	if(rvalid) if(is_last) num_chunk_elements = _IntNarrow_5_out;
	if(rvalid) if(!is_last) num_chunk_elements = _87;
end
always_comb begin // combinatorial is_last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_last = 1'bx;
	if(rvalid) is_last = _81;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_last = is_last;
end
always_comb begin // combinatorial _IntNarrow_5_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_5_in = 3'sdx;
	if(rvalid) if(is_last) _IntNarrow_5_in = _85;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _99;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial chunk_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_addr = 61'dx;
	if(request_new_burst) chunk_addr = _BitwiseIntSplit_2_upper;
end
always_comb begin // combinatorial element_in_chunk_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_in_chunk_align = 1'dx;
	if(request_new_burst) element_in_chunk_align = _BitwiseIntSplit_2_lower;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	element_in_chunk_align = element_in_chunk_align;
end
always_comb begin // combinatorial _BitwiseIntSplit_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_2_v = 62'dx;
	if(request_new_burst) _BitwiseIntSplit_2_v = _101;
end
always_comb begin // combinatorial chunk_count_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_count_bits = 33'dx;
	if(request_new_burst) chunk_count_bits = _BitwiseIntSplit_3_upper;
end
always_comb begin // combinatorial final_alignment
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	final_alignment = 1'dx;
	if(request_new_burst) final_alignment = _BitwiseIntSplit_3_lower;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	final_alignment = final_alignment;
end
always_comb begin // combinatorial _BitwiseIntSplit_3_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_3_v = 34'dx;
	if(request_new_burst) _BitwiseIntSplit_3_v = _104;
end
always_comb begin // combinatorial num_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunks = 33'dx;
	if(request_new_burst) if(is_no_chunks) num_chunks = 1'd1;
	if(request_new_burst) if(!is_no_chunks) num_chunks = _114;
end
always_comb begin // combinatorial is_no_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_no_chunks = 1'bx;
	if(request_new_burst) is_no_chunks = _107;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_no_chunks = is_no_chunks;
end
always_comb begin // combinatorial _BoolToInt_2_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_2_i = 1'bx;
	if(request_new_burst) if(!is_no_chunks) _BoolToInt_2_i = _113;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_2_i = _BoolToInt_2_i;
end
always_comb begin // combinatorial _BoolToInt_3_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_3_i = 1'bx;
	if(request_new_burst) _BoolToInt_3_i = _124;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_3_i = _BoolToInt_3_i;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_upper = 1'dx;
	if(request_new_burst) _BitwiseIntConcat_3_upper = _BoolToInt_3_o;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BitwiseIntConcat_3_upper = _BitwiseIntConcat_3_upper;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_lower = 1'dx;
	if(request_new_burst) _BitwiseIntConcat_3_lower = final_alignment;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BitwiseIntConcat_3_lower = _BitwiseIntConcat_3_lower;
end
always_comb begin // combinatorial _cur_start_chunk_addr_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_rst = 1'bx;
	_cur_start_chunk_addr_rst = _128;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_rst = _cur_start_chunk_addr_rst;
end
always_comb begin // combinatorial _num_chunks_left_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_rst = 1'bx;
	_num_chunks_left_rst = _130;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_rst = _num_chunks_left_rst;
end
endmodule

// BitwiseIntConcat #(UPPER_TO: 2, LOWER_BITS: 1)
module BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_1(
	input clk,
	input wire[0:0] upper,
	input wire[0:0] lower,
	output /*mux_wire*/ logic[1:0] v
);

/*mux_wire*/ logic[1:0] v_bits;
/*mux_wire*/ logic[0:0] _UIntToBits_value;
wire[0:0] _UIntToBits_bits;
/*mux_wire*/ logic[0:0] _UIntToBits_2_value;
wire[0:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[1:0] _FromBits_bits;
wire[1:0] _FromBits_value;
UIntToBits_NUM_BITS_1 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_1 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_4 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 2'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 2'bxx;
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
v_bits[1 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 1'dx;
	_UIntToBits_value = lower;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_UIntToBits_value = _UIntToBits_value;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 1'dx;
	_UIntToBits_2_value = upper;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_UIntToBits_2_value = _UIntToBits_2_value;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 2'bxx;
	_FromBits_bits = v_bits;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 4))
module FromBits_T_type_int_FROM_0_TO_4(
	input clk,
	input wire[1:0] bits,
	output /*mux_wire*/ logic[1:0] value
);

assign value = bits;
endmodule

// BitwiseIntSplit #(TO: 8589934593, LOWER_BITS: 1)
module BitwiseIntSplit_TO_8589934593_LOWER_BITS_1(
	input clk,
	input wire[33:0] v,
	output /*mux_wire*/ logic[32:0] upper,
	output /*mux_wire*/ logic[0:0] lower
);

genvar _g0;
/*mux_wire*/ logic[33:0] v_bits;
/*mux_wire*/ logic[33:0] _UIntToBits_value;
wire[33:0] _UIntToBits_bits;
wire[0:0] _2;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[0:0] _BitsToUInt_bits;
wire[0:0] _BitsToUInt_value;
wire[32:0] _3;
generate
for(_g0 = 0; _g0 < 33; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[1 + _g0];
end
endgenerate
/*mux_wire*/ logic[32:0] _FromBits_bits;
wire[32:0] _FromBits_value;
UIntToBits_NUM_BITS_34 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_1 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_4294967297 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 33'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 1'dx;
	lower = _BitsToUInt_value;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	lower = lower;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 34'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 34'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 1'bx;
	_BitsToUInt_bits = _2;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BitsToUInt_bits = _BitsToUInt_bits;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 4294967297))
module FromBits_T_type_int_FROM_0_TO_4294967297(
	input clk,
	input wire[32:0] bits,
	output /*mux_wire*/ logic[32:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 34)
module UIntToBits_NUM_BITS_34(
	input clk,
	input wire[33:0] value,
	output /*mux_wire*/ logic[33:0] bits
);

	assign bits = value;
endmodule

// BitwiseIntSplit #(TO: 4611686018427387904, LOWER_BITS: 1)
module BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_1(
	input clk,
	input wire[61:0] v,
	output /*mux_wire*/ logic[60:0] upper,
	output /*mux_wire*/ logic[0:0] lower
);

genvar _g0;
/*mux_wire*/ logic[61:0] v_bits;
/*mux_wire*/ logic[61:0] _UIntToBits_value;
wire[61:0] _UIntToBits_bits;
wire[0:0] _2;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[0:0] _BitsToUInt_bits;
wire[0:0] _BitsToUInt_value;
wire[60:0] _3;
generate
for(_g0 = 0; _g0 < 61; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[1 + _g0];
end
endgenerate
/*mux_wire*/ logic[60:0] _FromBits_bits;
wire[60:0] _FromBits_value;
UIntToBits_NUM_BITS_62 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_1 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_2305843009213693952 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 61'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 1'dx;
	lower = _BitsToUInt_value;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	lower = lower;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 62'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 62'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 1'bx;
	_BitsToUInt_bits = _2;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BitsToUInt_bits = _BitsToUInt_bits;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 61'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// BitsToUInt #(NUM_BITS: 1)
module BitsToUInt_NUM_BITS_1(
	input clk,
	input wire[0:0] bits,
	output /*mux_wire*/ logic[0:0] value
);

	assign value = bits;
endmodule

// IntNarrow #(FROM_I: -1, TO_I: 4, FROM: 0, TO: 3)
module IntNarrow_FROM_I_1_TO_I_4_FROM_0_TO_3(
	input clk,
	input wire signed[2:0] in,
	output /*mux_wire*/ logic[1:0] out
);

	assign out = in;
endmodule

// benchmark_burst_read #(AXI_WIDTH: 32)
module benchmark_burst_read_AXI_WIDTH_32(
	input aclk,
	input wire aresetn,
	input wire[11:0] s_axi_control_awaddr,
	input wire s_axi_control_awvalid,
	output /*mux_wire*/ logic s_axi_control_awready,
	input wire[31:0] s_axi_control_wdata,
	input wire[3:0] s_axi_control_wstrb,
	input wire s_axi_control_wvalid,
	output /*mux_wire*/ logic s_axi_control_wready,
	output /*mux_wire*/ logic[1:0] s_axi_control_bresp,
	output /*mux_wire*/ logic s_axi_control_bvalid,
	input wire s_axi_control_bready,
	input wire[11:0] s_axi_control_araddr,
	input wire s_axi_control_arvalid,
	output /*mux_wire*/ logic s_axi_control_arready,
	output /*mux_wire*/ logic[31:0] s_axi_control_rdata,
	output /*mux_wire*/ logic[1:0] s_axi_control_rresp,
	output /*mux_wire*/ logic s_axi_control_rvalid,
	input wire s_axi_control_rready,
	output /*mux_wire*/ logic m_axi_awvalid,
	input wire m_axi_awready,
	output /*mux_wire*/ logic[63:0] m_axi_awaddr,
	output /*mux_wire*/ logic[7:0] m_axi_awlen,
	output /*mux_wire*/ logic[1:0] m_axi_awburst,
	output /*mux_wire*/ logic[3:0] m_axi_awcache,
	output /*mux_wire*/ logic m_axi_wvalid,
	input wire m_axi_wready,
	output /*mux_wire*/ logic[31:0] m_axi_wdata,
	output /*mux_wire*/ logic[3:0] m_axi_wstrb,
	output /*mux_wire*/ logic m_axi_wlast,
	input wire m_axi_bvalid,
	output /*mux_wire*/ logic m_axi_bready,
	input wire[1:0] m_axi_bresp,
	output /*mux_wire*/ logic m_axi_arvalid,
	input wire m_axi_arready,
	output /*mux_wire*/ logic[63:0] m_axi_araddr,
	output /*mux_wire*/ logic[7:0] m_axi_arlen,
	output /*mux_wire*/ logic[2:0] m_axi_arsize,
	output /*mux_wire*/ logic[1:0] m_axi_arburst,
	input wire m_axi_rvalid,
	output /*mux_wire*/ logic m_axi_rready,
	input wire[31:0] m_axi_rdata,
	input wire[1:0] m_axi_rresp,
	input wire m_axi_rlast,
	output /*mux_wire*/ logic[2:0] m_axi_arprot,
	output /*mux_wire*/ logic[3:0] m_axi_arcache,
	output /*mux_wire*/ logic[3:0] m_axi_arqos,
	output /*mux_wire*/ logic m_axi_arlock,
	output /*mux_wire*/ logic[3:0] m_axi_arregion
);

genvar _g0;
/*mux_wire*/ logic _ctrl_aresetn;
wire _ctrl_awready;
wire _ctrl_wready;
wire[1:0] _ctrl_bresp;
wire _ctrl_bvalid;
wire _ctrl_arready;
wire[31:0] _ctrl_rdata;
wire[1:0] _ctrl_rresp;
wire _ctrl_rvalid;
/*mux_wire*/ logic[11:0] _ctrl_awaddr;
/*mux_wire*/ logic _ctrl_awvalid;
/*mux_wire*/ logic[31:0] _ctrl_wdata;
/*mux_wire*/ logic[3:0] _ctrl_wstrb;
/*mux_wire*/ logic _ctrl_wvalid;
/*mux_wire*/ logic _ctrl_bready;
/*mux_wire*/ logic[11:0] _ctrl_araddr;
/*mux_wire*/ logic _ctrl_arvalid;
/*mux_wire*/ logic _ctrl_rready;
/*mux_wire*/ logic _reader_aresetn;
/*mux_wire*/ logic _writer_aresetn;
wire _writer_awvalid;
wire[63:0] _writer_awaddr;
wire[7:0] _writer_awlen;
wire[1:0] _writer_awburst;
wire[3:0] _writer_awcache;
wire _writer_wvalid;
wire[31:0] _writer_wdata;
wire[3:0] _writer_wstrb;
wire _writer_wlast;
wire _writer_bready;
/*mux_wire*/ logic _writer_awready;
/*mux_wire*/ logic _writer_wready;
/*mux_wire*/ logic _writer_bvalid;
/*mux_wire*/ logic[1:0] _writer_bresp;
wire _reader_arvalid;
wire[63:0] _reader_araddr;
wire[7:0] _reader_arlen;
wire[2:0] _reader_arsize;
wire[1:0] _reader_arburst;
wire _reader_rready;
/*mux_wire*/ logic _reader_arready;
/*mux_wire*/ logic _reader_rvalid;
/*mux_wire*/ logic[31:0] _reader_rdata;
/*mux_wire*/ logic[1:0] _reader_rresp;
/*mux_wire*/ logic _reader_rlast;
/*mux_wire*/ logic[63:0] addr_a_bits;
wire[31:0] _ctrl_input_regs[3:0];
wire[31:0] _46 = _ctrl_input_regs[0];
wire[31:0] _47 = _ctrl_input_regs[1];
/*mux_wire*/ logic[63:0] start_addr;
/*mux_wire*/ logic[63:0] _BitsToUInt_bits;
wire[63:0] _BitsToUInt_value;
/*mux_wire*/ logic[31:0] num_to_transfer;
wire[31:0] _49 = _ctrl_input_regs[2];
/*mux_wire*/ logic[31:0] _BitsToUInt_2_bits;
wire[31:0] _BitsToUInt_2_value;
/*mux_wire*/ logic[31:0] _IntNarrow_in;
wire[31:0] _IntNarrow_out;
/*mux_wire*/ logic[31:0] config_bits;
wire[31:0] _50 = _ctrl_input_regs[3];
wire[2:0] _51;
generate
for(_g0 = 0; _g0 < 3; _g0 = _g0 + 1) begin
assign _51[_g0] = config_bits[5 + _g0];
end
endgenerate
wire[3:0] _52;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _52[_g0] = config_bits[8 + _g0];
end
endgenerate
wire[3:0] _53;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _53[_g0] = config_bits[12 + _g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_3_bits;
wire[3:0] _BitsToUInt_3_value;
wire _54 = config_bits[16];
wire[3:0] _55;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _55[_g0] = config_bits[17 + _g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_4_bits;
wire[3:0] _BitsToUInt_4_value;
wire[10:0] _56;
generate
for(_g0 = 0; _g0 < 11; _g0 = _g0 + 1) begin
assign _56[_g0] = config_bits[21 + _g0];
end
endgenerate
/*mux_wire*/ logic[10:0] _BitsToUInt_5_bits;
wire[10:0] _BitsToUInt_5_value;
/*mux_wire*/ logic[10:0] _reader_max_in_flight;
/*state*/ logic[63:0] cycles_since_reset;
wire[64:0] _59;
assign _59 = cycles_since_reset + 1'd1;
wire[63:0] _60;
assign _60 = _59; // == mod 18446744073709551616 (target is 64 bits wide)
/*mux_wire*/ logic[63:0] cycles_since_reset_bits;
/*mux_wire*/ logic[63:0] _UIntToBits_value;
wire[63:0] _UIntToBits_bits;
/*latency*/ logic[63:0] __UIntToBits_bits_D1; always_ff @(posedge aclk) begin __UIntToBits_bits_D1 <= _UIntToBits_bits; end
/*latency*/ logic[63:0] __UIntToBits_bits_D2; always_ff @(posedge aclk) begin __UIntToBits_bits_D2 <= __UIntToBits_bits_D1; end
/*latency*/ logic[63:0] __UIntToBits_bits_D3; always_ff @(posedge aclk) begin __UIntToBits_bits_D3 <= __UIntToBits_bits_D2; end
/*state*/ logic[63:0] cycles_since_reset_at_start;
/*state*/ logic running;
/*state*/ logic[31:0] num_cycles_running;
/*state*/ logic[31:0] hash;
wire _ctrl_start;
/*latency*/ logic __ctrl_start_D1; always_ff @(posedge aclk) begin __ctrl_start_D1 <= _ctrl_start; end
/*latency*/ logic __ctrl_start_D2; always_ff @(posedge aclk) begin __ctrl_start_D2 <= __ctrl_start_D1; end
/*latency*/ logic __ctrl_start_D3; always_ff @(posedge aclk) begin __ctrl_start_D3 <= __ctrl_start_D2; end
/*mux_wire*/ logic _reader_request_new_burst;
/*mux_wire*/ logic[63:0] _reader_start_addr;
/*mux_wire*/ logic[31:0] _reader_count;
localparam[31:0] _67 = 32'b00000000000000000000000000000000;
wire[32:0] _72;
assign _72 = num_cycles_running + 1'd1;
wire[31:0] _73;
assign _73 = _72; // == mod 4294967296 (target is 32 bits wide)
/*mux_wire*/ logic _reader_is_ready_to_receive_lots_of_data;
wire _reader_value_valid;
/*latency*/ logic __reader_value_valid_D1; always_ff @(posedge aclk) begin __reader_value_valid_D1 <= _reader_value_valid; end
/*latency*/ logic __reader_value_valid_D2; always_ff @(posedge aclk) begin __reader_value_valid_D2 <= __reader_value_valid_D1; end
/*latency*/ logic __reader_value_valid_D3; always_ff @(posedge aclk) begin __reader_value_valid_D3 <= __reader_value_valid_D2; end
wire[31:0] _reader_value[0:0];
wire _reader_last;
/*mux_wire*/ logic[31:0] value[0:0];
/*mux_wire*/ logic last;
/*latency*/ logic _last_D1; always_ff @(posedge aclk) begin _last_D1 <= last; end
/*latency*/ logic _last_D2; always_ff @(posedge aclk) begin _last_D2 <= _last_D1; end
/*latency*/ logic _last_D3; always_ff @(posedge aclk) begin _last_D3 <= _last_D2; end
/*mux_wire*/ logic[31:0] new_hash_contrib;
wire[0:0] _74;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _74[_g0] = value[_g0][0];
end
endgenerate
wire _75;
assign _75 = ^_74;
/*latency*/ logic __75_D1; always_ff @(posedge aclk) begin __75_D1 <= _75; end
/*latency*/ logic __75_D2; always_ff @(posedge aclk) begin __75_D2 <= __75_D1; end
wire[0:0] _76;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _76[_g0] = value[_g0][1];
end
endgenerate
wire _77;
assign _77 = ^_76;
/*latency*/ logic __77_D1; always_ff @(posedge aclk) begin __77_D1 <= _77; end
/*latency*/ logic __77_D2; always_ff @(posedge aclk) begin __77_D2 <= __77_D1; end
wire[0:0] _78;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _78[_g0] = value[_g0][2];
end
endgenerate
wire _79;
assign _79 = ^_78;
/*latency*/ logic __79_D1; always_ff @(posedge aclk) begin __79_D1 <= _79; end
/*latency*/ logic __79_D2; always_ff @(posedge aclk) begin __79_D2 <= __79_D1; end
wire[0:0] _80;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _80[_g0] = value[_g0][3];
end
endgenerate
wire _81;
assign _81 = ^_80;
/*latency*/ logic __81_D1; always_ff @(posedge aclk) begin __81_D1 <= _81; end
/*latency*/ logic __81_D2; always_ff @(posedge aclk) begin __81_D2 <= __81_D1; end
wire[0:0] _82;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _82[_g0] = value[_g0][4];
end
endgenerate
wire _83;
assign _83 = ^_82;
/*latency*/ logic __83_D1; always_ff @(posedge aclk) begin __83_D1 <= _83; end
/*latency*/ logic __83_D2; always_ff @(posedge aclk) begin __83_D2 <= __83_D1; end
wire[0:0] _84;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _84[_g0] = value[_g0][5];
end
endgenerate
wire _85;
assign _85 = ^_84;
/*latency*/ logic __85_D1; always_ff @(posedge aclk) begin __85_D1 <= _85; end
/*latency*/ logic __85_D2; always_ff @(posedge aclk) begin __85_D2 <= __85_D1; end
wire[0:0] _86;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _86[_g0] = value[_g0][6];
end
endgenerate
wire _87;
assign _87 = ^_86;
/*latency*/ logic __87_D1; always_ff @(posedge aclk) begin __87_D1 <= _87; end
/*latency*/ logic __87_D2; always_ff @(posedge aclk) begin __87_D2 <= __87_D1; end
wire[0:0] _88;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _88[_g0] = value[_g0][7];
end
endgenerate
wire _89;
assign _89 = ^_88;
/*latency*/ logic __89_D1; always_ff @(posedge aclk) begin __89_D1 <= _89; end
/*latency*/ logic __89_D2; always_ff @(posedge aclk) begin __89_D2 <= __89_D1; end
wire[0:0] _90;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _90[_g0] = value[_g0][8];
end
endgenerate
wire _91;
assign _91 = ^_90;
/*latency*/ logic __91_D1; always_ff @(posedge aclk) begin __91_D1 <= _91; end
/*latency*/ logic __91_D2; always_ff @(posedge aclk) begin __91_D2 <= __91_D1; end
wire[0:0] _92;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _92[_g0] = value[_g0][9];
end
endgenerate
wire _93;
assign _93 = ^_92;
/*latency*/ logic __93_D1; always_ff @(posedge aclk) begin __93_D1 <= _93; end
/*latency*/ logic __93_D2; always_ff @(posedge aclk) begin __93_D2 <= __93_D1; end
wire[0:0] _94;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _94[_g0] = value[_g0][10];
end
endgenerate
wire _95;
assign _95 = ^_94;
/*latency*/ logic __95_D1; always_ff @(posedge aclk) begin __95_D1 <= _95; end
/*latency*/ logic __95_D2; always_ff @(posedge aclk) begin __95_D2 <= __95_D1; end
wire[0:0] _96;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _96[_g0] = value[_g0][11];
end
endgenerate
wire _97;
assign _97 = ^_96;
/*latency*/ logic __97_D1; always_ff @(posedge aclk) begin __97_D1 <= _97; end
/*latency*/ logic __97_D2; always_ff @(posedge aclk) begin __97_D2 <= __97_D1; end
wire[0:0] _98;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _98[_g0] = value[_g0][12];
end
endgenerate
wire _99;
assign _99 = ^_98;
/*latency*/ logic __99_D1; always_ff @(posedge aclk) begin __99_D1 <= _99; end
/*latency*/ logic __99_D2; always_ff @(posedge aclk) begin __99_D2 <= __99_D1; end
wire[0:0] _100;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _100[_g0] = value[_g0][13];
end
endgenerate
wire _101;
assign _101 = ^_100;
/*latency*/ logic __101_D1; always_ff @(posedge aclk) begin __101_D1 <= _101; end
/*latency*/ logic __101_D2; always_ff @(posedge aclk) begin __101_D2 <= __101_D1; end
wire[0:0] _102;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _102[_g0] = value[_g0][14];
end
endgenerate
wire _103;
assign _103 = ^_102;
/*latency*/ logic __103_D1; always_ff @(posedge aclk) begin __103_D1 <= _103; end
/*latency*/ logic __103_D2; always_ff @(posedge aclk) begin __103_D2 <= __103_D1; end
wire[0:0] _104;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _104[_g0] = value[_g0][15];
end
endgenerate
wire _105;
assign _105 = ^_104;
/*latency*/ logic __105_D1; always_ff @(posedge aclk) begin __105_D1 <= _105; end
/*latency*/ logic __105_D2; always_ff @(posedge aclk) begin __105_D2 <= __105_D1; end
wire[0:0] _106;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _106[_g0] = value[_g0][16];
end
endgenerate
wire _107;
assign _107 = ^_106;
/*latency*/ logic __107_D1; always_ff @(posedge aclk) begin __107_D1 <= _107; end
/*latency*/ logic __107_D2; always_ff @(posedge aclk) begin __107_D2 <= __107_D1; end
wire[0:0] _108;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _108[_g0] = value[_g0][17];
end
endgenerate
wire _109;
assign _109 = ^_108;
/*latency*/ logic __109_D1; always_ff @(posedge aclk) begin __109_D1 <= _109; end
/*latency*/ logic __109_D2; always_ff @(posedge aclk) begin __109_D2 <= __109_D1; end
wire[0:0] _110;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _110[_g0] = value[_g0][18];
end
endgenerate
wire _111;
assign _111 = ^_110;
/*latency*/ logic __111_D1; always_ff @(posedge aclk) begin __111_D1 <= _111; end
/*latency*/ logic __111_D2; always_ff @(posedge aclk) begin __111_D2 <= __111_D1; end
wire[0:0] _112;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _112[_g0] = value[_g0][19];
end
endgenerate
wire _113;
assign _113 = ^_112;
/*latency*/ logic __113_D1; always_ff @(posedge aclk) begin __113_D1 <= _113; end
/*latency*/ logic __113_D2; always_ff @(posedge aclk) begin __113_D2 <= __113_D1; end
wire[0:0] _114;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _114[_g0] = value[_g0][20];
end
endgenerate
wire _115;
assign _115 = ^_114;
/*latency*/ logic __115_D1; always_ff @(posedge aclk) begin __115_D1 <= _115; end
/*latency*/ logic __115_D2; always_ff @(posedge aclk) begin __115_D2 <= __115_D1; end
wire[0:0] _116;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _116[_g0] = value[_g0][21];
end
endgenerate
wire _117;
assign _117 = ^_116;
/*latency*/ logic __117_D1; always_ff @(posedge aclk) begin __117_D1 <= _117; end
/*latency*/ logic __117_D2; always_ff @(posedge aclk) begin __117_D2 <= __117_D1; end
wire[0:0] _118;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _118[_g0] = value[_g0][22];
end
endgenerate
wire _119;
assign _119 = ^_118;
/*latency*/ logic __119_D1; always_ff @(posedge aclk) begin __119_D1 <= _119; end
/*latency*/ logic __119_D2; always_ff @(posedge aclk) begin __119_D2 <= __119_D1; end
wire[0:0] _120;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _120[_g0] = value[_g0][23];
end
endgenerate
wire _121;
assign _121 = ^_120;
/*latency*/ logic __121_D1; always_ff @(posedge aclk) begin __121_D1 <= _121; end
/*latency*/ logic __121_D2; always_ff @(posedge aclk) begin __121_D2 <= __121_D1; end
wire[0:0] _122;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _122[_g0] = value[_g0][24];
end
endgenerate
wire _123;
assign _123 = ^_122;
/*latency*/ logic __123_D1; always_ff @(posedge aclk) begin __123_D1 <= _123; end
/*latency*/ logic __123_D2; always_ff @(posedge aclk) begin __123_D2 <= __123_D1; end
wire[0:0] _124;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _124[_g0] = value[_g0][25];
end
endgenerate
wire _125;
assign _125 = ^_124;
/*latency*/ logic __125_D1; always_ff @(posedge aclk) begin __125_D1 <= _125; end
/*latency*/ logic __125_D2; always_ff @(posedge aclk) begin __125_D2 <= __125_D1; end
wire[0:0] _126;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _126[_g0] = value[_g0][26];
end
endgenerate
wire _127;
assign _127 = ^_126;
/*latency*/ logic __127_D1; always_ff @(posedge aclk) begin __127_D1 <= _127; end
/*latency*/ logic __127_D2; always_ff @(posedge aclk) begin __127_D2 <= __127_D1; end
wire[0:0] _128;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _128[_g0] = value[_g0][27];
end
endgenerate
wire _129;
assign _129 = ^_128;
/*latency*/ logic __129_D1; always_ff @(posedge aclk) begin __129_D1 <= _129; end
/*latency*/ logic __129_D2; always_ff @(posedge aclk) begin __129_D2 <= __129_D1; end
wire[0:0] _130;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _130[_g0] = value[_g0][28];
end
endgenerate
wire _131;
assign _131 = ^_130;
/*latency*/ logic __131_D1; always_ff @(posedge aclk) begin __131_D1 <= _131; end
/*latency*/ logic __131_D2; always_ff @(posedge aclk) begin __131_D2 <= __131_D1; end
wire[0:0] _132;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _132[_g0] = value[_g0][29];
end
endgenerate
wire _133;
assign _133 = ^_132;
/*latency*/ logic __133_D1; always_ff @(posedge aclk) begin __133_D1 <= _133; end
/*latency*/ logic __133_D2; always_ff @(posedge aclk) begin __133_D2 <= __133_D1; end
wire[0:0] _134;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _134[_g0] = value[_g0][30];
end
endgenerate
wire _135;
assign _135 = ^_134;
/*latency*/ logic __135_D1; always_ff @(posedge aclk) begin __135_D1 <= _135; end
/*latency*/ logic __135_D2; always_ff @(posedge aclk) begin __135_D2 <= __135_D1; end
wire[0:0] _136;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _136[_g0] = value[_g0][31];
end
endgenerate
wire _137;
assign _137 = ^_136;
/*latency*/ logic __137_D1; always_ff @(posedge aclk) begin __137_D1 <= _137; end
/*latency*/ logic __137_D2; always_ff @(posedge aclk) begin __137_D2 <= __137_D1; end
/*mux_wire*/ logic[31:0] new_hash;
/*latency*/ logic[31:0] _new_hash_D3; always_ff @(posedge aclk) begin _new_hash_D3 <= new_hash; end
wire[31:0] _140;
assign _140 = hash ^ new_hash_contrib;
/*mux_wire*/ logic[31:0] _UIntToBits_2_value;
wire[31:0] _UIntToBits_2_bits;
/*latency*/ logic[31:0] __UIntToBits_2_bits_D1; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D1 <= _UIntToBits_2_bits; end
/*latency*/ logic[31:0] __UIntToBits_2_bits_D2; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D2 <= __UIntToBits_2_bits_D1; end
/*latency*/ logic[31:0] __UIntToBits_2_bits_D3; always_ff @(posedge aclk) begin __UIntToBits_2_bits_D3 <= __UIntToBits_2_bits_D2; end
wire[31:0] _144;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _144[_g0] = cycles_since_reset_at_start[_g0];
end
endgenerate
wire[31:0] _145;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _145[_g0] = cycles_since_reset_at_start[32 + _g0];
end
endgenerate
wire[31:0] _146;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _146[_g0] = cycles_since_reset_bits[_g0];
end
endgenerate
wire[31:0] _147;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _147[_g0] = cycles_since_reset_bits[32 + _g0];
end
endgenerate
wire[31:0] _148[5:0];
assign _148[0] = __UIntToBits_2_bits_D3;
assign _148[1] = _new_hash_D3;
assign _148[2] = _144;
assign _148[3] = _145;
assign _148[4] = _146;
assign _148[5] = _147;
/*mux_wire*/ logic _ctrl_finish;
/*mux_wire*/ logic[31:0] _ctrl_output_regs[5:0];
wire _153;
assign _153 = !aresetn;
/*latency*/ logic __153_D1; always_ff @(posedge aclk) begin __153_D1 <= _153; end
/*latency*/ logic __153_D2; always_ff @(posedge aclk) begin __153_D2 <= __153_D1; end
localparam[31:0] _155 = 32'b00000000000000000000000000000000;
axi_ctrl_slave_NUM_INPUT_REGS_4_NUM_OUTPUT_REGS_6_ADDR_WIDTH_12_AXI_WIDTH_32 ctrl(
	.aclk(aclk),
	.aresetn(_ctrl_aresetn),
	.awaddr(_ctrl_awaddr),
	.awvalid(_ctrl_awvalid),
	.awready(_ctrl_awready),
	.wdata(_ctrl_wdata),
	.wstrb(_ctrl_wstrb),
	.wvalid(_ctrl_wvalid),
	.wready(_ctrl_wready),
	.bresp(_ctrl_bresp),
	.bvalid(_ctrl_bvalid),
	.bready(_ctrl_bready),
	.araddr(_ctrl_araddr),
	.arvalid(_ctrl_arvalid),
	.arready(_ctrl_arready),
	.rdata(_ctrl_rdata),
	.rresp(_ctrl_rresp),
	.rvalid(_ctrl_rvalid),
	.rready(_ctrl_rready),
	.input_regs(_ctrl_input_regs),
	.start(_ctrl_start),
	.finish(_ctrl_finish),
	.output_regs(_ctrl_output_regs)
);
axi_realigning_burst_reader_T_type_bool_32_1_AXI_WIDTH_32_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616 reader(
	.aclk(aclk),
	.aresetn(_reader_aresetn),
	.arvalid(_reader_arvalid),
	.arready(_reader_arready),
	.araddr(_reader_araddr),
	.arlen(_reader_arlen),
	.arsize(_reader_arsize),
	.arburst(_reader_arburst),
	.arprot(),
	.arcache(),
	.arqos(),
	.arlock(),
	.arregion(),
	.rvalid(_reader_rvalid),
	.rready(_reader_rready),
	.rdata(_reader_rdata),
	.rresp(_reader_rresp),
	.rlast(_reader_rlast),
	.max_in_flight(_reader_max_in_flight),
	.may_request_new_burst(),
	.request_new_burst(_reader_request_new_burst),
	.start_addr(_reader_start_addr),
	.count(_reader_count),
	.is_ready_to_receive_lots_of_data(_reader_is_ready_to_receive_lots_of_data),
	.value_valid(_reader_value_valid),
	.value(_reader_value),
	.last(_reader_last)
);
axi_memory_writer_tie_off_AXI_WIDTH_32 writer(
	.aclk(aclk),
	.aresetn(_writer_aresetn),
	.awvalid(_writer_awvalid),
	.awready(_writer_awready),
	.awaddr(_writer_awaddr),
	.awlen(_writer_awlen),
	.awsize(),
	.awburst(_writer_awburst),
	.awprot(),
	.awcache(_writer_awcache),
	.awqos(),
	.awlock(),
	.awregion(),
	.wvalid(_writer_wvalid),
	.wready(_writer_wready),
	.wdata(_writer_wdata),
	.wstrb(_writer_wstrb),
	.wlast(_writer_wlast),
	.bvalid(_writer_bvalid),
	.bresp(_writer_bresp),
	.bready(_writer_bready)
);
BitsToUInt_NUM_BITS_64 BitsToUInt(
	.clk(aclk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
BitsToUInt_NUM_BITS_32 BitsToUInt_2(
	.clk(aclk),
	.bits(_BitsToUInt_2_bits),
	.value(_BitsToUInt_2_value)
);
IntNarrow_FROM_I_0_TO_I_4294967296_FROM_1_TO_4294967296 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
BitsToUInt_NUM_BITS_4 BitsToUInt_3(
	.clk(aclk),
	.bits(_BitsToUInt_3_bits),
	.value(_BitsToUInt_3_value)
);
BitsToUInt_NUM_BITS_4 BitsToUInt_4(
	.clk(aclk),
	.bits(_BitsToUInt_4_bits),
	.value(_BitsToUInt_4_value)
);
BitsToUInt_NUM_BITS_11 BitsToUInt_5(
	.clk(aclk),
	.bits(_BitsToUInt_5_bits),
	.value(_BitsToUInt_5_value)
);
UIntToBits_NUM_BITS_64 UIntToBits(
	.clk(aclk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_32 UIntToBits_2(
	.clk(aclk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
always_comb begin // combinatorial _ctrl_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_aresetn = 1'bx;
	_ctrl_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_aresetn = _ctrl_aresetn;
end
always_comb begin // combinatorial s_axi_control_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_awready = 1'bx;
	s_axi_control_awready = _ctrl_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_awready = s_axi_control_awready;
end
always_comb begin // combinatorial s_axi_control_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_wready = 1'bx;
	s_axi_control_wready = _ctrl_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_wready = s_axi_control_wready;
end
always_comb begin // combinatorial s_axi_control_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bresp = 2'bxx;
	s_axi_control_bresp = _ctrl_bresp;
end
always_comb begin // combinatorial s_axi_control_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bvalid = 1'bx;
	s_axi_control_bvalid = _ctrl_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_bvalid = s_axi_control_bvalid;
end
always_comb begin // combinatorial s_axi_control_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_arready = 1'bx;
	s_axi_control_arready = _ctrl_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_arready = s_axi_control_arready;
end
always_comb begin // combinatorial s_axi_control_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	s_axi_control_rdata = _ctrl_rdata;
end
always_comb begin // combinatorial s_axi_control_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rresp = 2'bxx;
	s_axi_control_rresp = _ctrl_rresp;
end
always_comb begin // combinatorial s_axi_control_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rvalid = 1'bx;
	s_axi_control_rvalid = _ctrl_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_rvalid = s_axi_control_rvalid;
end
always_comb begin // combinatorial _ctrl_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awaddr = 12'dx;
	_ctrl_awaddr = s_axi_control_awaddr;
end
always_comb begin // combinatorial _ctrl_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awvalid = 1'bx;
	_ctrl_awvalid = s_axi_control_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_awvalid = _ctrl_awvalid;
end
always_comb begin // combinatorial _ctrl_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_ctrl_wdata = s_axi_control_wdata;
end
always_comb begin // combinatorial _ctrl_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wstrb = 4'bxxxx;
	_ctrl_wstrb = s_axi_control_wstrb;
end
always_comb begin // combinatorial _ctrl_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wvalid = 1'bx;
	_ctrl_wvalid = s_axi_control_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_wvalid = _ctrl_wvalid;
end
always_comb begin // combinatorial _ctrl_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_bready = 1'bx;
	_ctrl_bready = s_axi_control_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_bready = _ctrl_bready;
end
always_comb begin // combinatorial _ctrl_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_araddr = 12'dx;
	_ctrl_araddr = s_axi_control_araddr;
end
always_comb begin // combinatorial _ctrl_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_arvalid = 1'bx;
	_ctrl_arvalid = s_axi_control_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_arvalid = _ctrl_arvalid;
end
always_comb begin // combinatorial _ctrl_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_rready = 1'bx;
	_ctrl_rready = s_axi_control_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_rready = _ctrl_rready;
end
always_comb begin // combinatorial _reader_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_aresetn = 1'bx;
	_reader_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_aresetn = _reader_aresetn;
end
always_comb begin // combinatorial _writer_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_aresetn = 1'bx;
	_writer_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_aresetn = _writer_aresetn;
end
always_comb begin // combinatorial m_axi_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awvalid = 1'bx;
	m_axi_awvalid = _writer_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_awvalid = m_axi_awvalid;
end
always_comb begin // combinatorial m_axi_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awaddr = 64'dx;
	m_axi_awaddr = _writer_awaddr;
end
always_comb begin // combinatorial m_axi_awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awlen = 8'dx;
	m_axi_awlen = _writer_awlen;
end
always_comb begin // combinatorial m_axi_awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awburst = 2'bxx;
	m_axi_awburst = _writer_awburst;
end
always_comb begin // combinatorial m_axi_awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awcache = 4'bxxxx;
	m_axi_awcache = _writer_awcache;
end
always_comb begin // combinatorial m_axi_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wvalid = 1'bx;
	m_axi_wvalid = _writer_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wvalid = m_axi_wvalid;
end
always_comb begin // combinatorial m_axi_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	m_axi_wdata = _writer_wdata;
end
always_comb begin // combinatorial m_axi_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wstrb = 4'bxxxx;
	m_axi_wstrb = _writer_wstrb;
end
always_comb begin // combinatorial m_axi_wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wlast = 1'bx;
	m_axi_wlast = _writer_wlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wlast = m_axi_wlast;
end
always_comb begin // combinatorial m_axi_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_bready = 1'bx;
	m_axi_bready = _writer_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_bready = m_axi_bready;
end
always_comb begin // combinatorial _writer_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_awready = 1'bx;
	_writer_awready = m_axi_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_awready = _writer_awready;
end
always_comb begin // combinatorial _writer_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_wready = 1'bx;
	_writer_wready = m_axi_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_wready = _writer_wready;
end
always_comb begin // combinatorial _writer_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bvalid = 1'bx;
	_writer_bvalid = m_axi_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_bvalid = _writer_bvalid;
end
always_comb begin // combinatorial _writer_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bresp = 2'bxx;
	_writer_bresp = m_axi_bresp;
end
always_comb begin // combinatorial m_axi_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arvalid = 1'bx;
	m_axi_arvalid = _reader_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arvalid = m_axi_arvalid;
end
always_comb begin // combinatorial m_axi_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_araddr = 64'dx;
	m_axi_araddr = _reader_araddr;
end
always_comb begin // combinatorial m_axi_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlen = 8'dx;
	m_axi_arlen = _reader_arlen;
end
always_comb begin // combinatorial m_axi_arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arsize = 3'dx;
	m_axi_arsize = _reader_arsize;
end
always_comb begin // combinatorial m_axi_arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arburst = 2'bxx;
	m_axi_arburst = _reader_arburst;
end
always_comb begin // combinatorial m_axi_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_rready = 1'bx;
	m_axi_rready = _reader_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_rready = m_axi_rready;
end
always_comb begin // combinatorial _reader_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_arready = 1'bx;
	_reader_arready = m_axi_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_arready = _reader_arready;
end
always_comb begin // combinatorial _reader_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rvalid = 1'bx;
	_reader_rvalid = m_axi_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rvalid = _reader_rvalid;
end
always_comb begin // combinatorial _reader_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_reader_rdata = m_axi_rdata;
end
always_comb begin // combinatorial _reader_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rresp = 2'bxx;
	_reader_rresp = m_axi_rresp;
end
always_comb begin // combinatorial _reader_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rlast = 1'bx;
	_reader_rlast = m_axi_rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rlast = _reader_rlast;
end
always_comb begin // combinatorial addr_a_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	addr_a_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[_v0] = _46[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[32 + _v0] = _47[_v0];
end
end
always_comb begin // combinatorial start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	start_addr = 64'dx;
	start_addr = _BitsToUInt_value;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_BitsToUInt_bits = addr_a_bits;
end
always_comb begin // combinatorial num_to_transfer
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_to_transfer = 32'dx;
	num_to_transfer = _IntNarrow_out;
end
always_comb begin // combinatorial _BitsToUInt_2_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_2_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_BitsToUInt_2_bits = _49;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 32'dx;
	_IntNarrow_in = _BitsToUInt_2_value;
end
always_comb begin // combinatorial config_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	config_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	config_bits = _50;
end
always_comb begin // combinatorial m_axi_arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arprot = 3'bxxx;
	m_axi_arprot = _51;
end
always_comb begin // combinatorial m_axi_arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arcache = 4'bxxxx;
	m_axi_arcache = _52;
end
always_comb begin // combinatorial m_axi_arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arqos = 4'dx;
	m_axi_arqos = _BitsToUInt_3_value;
end
always_comb begin // combinatorial _BitsToUInt_3_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_3_bits = 4'bxxxx;
	_BitsToUInt_3_bits = _53;
end
always_comb begin // combinatorial m_axi_arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlock = 1'bx;
	m_axi_arlock = _54;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arlock = m_axi_arlock;
end
always_comb begin // combinatorial m_axi_arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arregion = 4'dx;
	m_axi_arregion = _BitsToUInt_4_value;
end
always_comb begin // combinatorial _BitsToUInt_4_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_4_bits = 4'bxxxx;
	_BitsToUInt_4_bits = _55;
end
always_comb begin // combinatorial _BitsToUInt_5_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_5_bits = 11'bxxxxxxxxxxx;
	_BitsToUInt_5_bits = _56;
end
always_comb begin // combinatorial _reader_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_max_in_flight = 11'dx;
	_reader_max_in_flight = _BitsToUInt_5_value;
end
always_ff @(posedge aclk) begin // state cycles_since_reset
	cycles_since_reset <= _60;
	if(_153) cycles_since_reset <= 1'd0;
end
always_comb begin // combinatorial cycles_since_reset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cycles_since_reset_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	cycles_since_reset_bits = __UIntToBits_bits_D3;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 64'dx;
	_UIntToBits_value = cycles_since_reset;
end
always_ff @(posedge aclk) begin // state cycles_since_reset_at_start
	if(__ctrl_start_D3) cycles_since_reset_at_start <= cycles_since_reset_bits;
end
always_ff @(posedge aclk) begin // state running
	if(_ctrl_start) running <= 1'b1;
	if(_reader_value_valid) if(last) running <= 1'b0;
	if(_153) running <= 1'b0;
end
always_ff @(posedge aclk) begin // state num_cycles_running
	if(_ctrl_start) num_cycles_running <= 1'd0;
	if(running) num_cycles_running <= _73;
	if(_153) num_cycles_running <= 1'd0;
end
always_ff @(posedge aclk) begin // state hash
	if(__ctrl_start_D2) hash <= _67;
	if(__reader_value_valid_D2) hash <= new_hash;
	if(__153_D2) hash <= _155;
end
always_comb begin // combinatorial _reader_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_request_new_burst = 1'bx;
	_reader_request_new_burst = 1'b0;
	if(_ctrl_start) _reader_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_request_new_burst = _reader_request_new_burst;
end
always_comb begin // combinatorial _reader_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_start_addr = 64'dx;
	if(_ctrl_start) _reader_start_addr = start_addr;
end
always_comb begin // combinatorial _reader_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_count = 32'dx;
	if(_ctrl_start) _reader_count = num_to_transfer;
end
always_comb begin // combinatorial _reader_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_is_ready_to_receive_lots_of_data = 1'bx;
	_reader_is_ready_to_receive_lots_of_data = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_is_ready_to_receive_lots_of_data = _reader_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_reader_value_valid) value[_v0] = _reader_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_reader_value_valid) last = _reader_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_comb begin // combinatorial new_hash_contrib
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_hash_contrib = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(__reader_value_valid_D2) new_hash_contrib[0] = __75_D2;
	if(__reader_value_valid_D2) new_hash_contrib[1] = __77_D2;
	if(__reader_value_valid_D2) new_hash_contrib[2] = __79_D2;
	if(__reader_value_valid_D2) new_hash_contrib[3] = __81_D2;
	if(__reader_value_valid_D2) new_hash_contrib[4] = __83_D2;
	if(__reader_value_valid_D2) new_hash_contrib[5] = __85_D2;
	if(__reader_value_valid_D2) new_hash_contrib[6] = __87_D2;
	if(__reader_value_valid_D2) new_hash_contrib[7] = __89_D2;
	if(__reader_value_valid_D2) new_hash_contrib[8] = __91_D2;
	if(__reader_value_valid_D2) new_hash_contrib[9] = __93_D2;
	if(__reader_value_valid_D2) new_hash_contrib[10] = __95_D2;
	if(__reader_value_valid_D2) new_hash_contrib[11] = __97_D2;
	if(__reader_value_valid_D2) new_hash_contrib[12] = __99_D2;
	if(__reader_value_valid_D2) new_hash_contrib[13] = __101_D2;
	if(__reader_value_valid_D2) new_hash_contrib[14] = __103_D2;
	if(__reader_value_valid_D2) new_hash_contrib[15] = __105_D2;
	if(__reader_value_valid_D2) new_hash_contrib[16] = __107_D2;
	if(__reader_value_valid_D2) new_hash_contrib[17] = __109_D2;
	if(__reader_value_valid_D2) new_hash_contrib[18] = __111_D2;
	if(__reader_value_valid_D2) new_hash_contrib[19] = __113_D2;
	if(__reader_value_valid_D2) new_hash_contrib[20] = __115_D2;
	if(__reader_value_valid_D2) new_hash_contrib[21] = __117_D2;
	if(__reader_value_valid_D2) new_hash_contrib[22] = __119_D2;
	if(__reader_value_valid_D2) new_hash_contrib[23] = __121_D2;
	if(__reader_value_valid_D2) new_hash_contrib[24] = __123_D2;
	if(__reader_value_valid_D2) new_hash_contrib[25] = __125_D2;
	if(__reader_value_valid_D2) new_hash_contrib[26] = __127_D2;
	if(__reader_value_valid_D2) new_hash_contrib[27] = __129_D2;
	if(__reader_value_valid_D2) new_hash_contrib[28] = __131_D2;
	if(__reader_value_valid_D2) new_hash_contrib[29] = __133_D2;
	if(__reader_value_valid_D2) new_hash_contrib[30] = __135_D2;
	if(__reader_value_valid_D2) new_hash_contrib[31] = __137_D2;
end
always_comb begin // combinatorial new_hash
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_hash = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(__reader_value_valid_D2) new_hash = _140;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 32'dx;
	if(_reader_value_valid) if(last) _UIntToBits_2_value = num_cycles_running;
end
always_comb begin // combinatorial _ctrl_finish
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_finish = 1'bx;
	_ctrl_finish = 1'b0;
	if(__reader_value_valid_D3) if(_last_D3) _ctrl_finish = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_finish = _ctrl_finish;
end
always_comb begin // combinatorial _ctrl_output_regs
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_output_regs = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
if(__reader_value_valid_D3) if(_last_D3) _ctrl_output_regs[_v0] = _148[_v0];
end
end
endmodule

// UIntToBits #(NUM_BITS: 64)
module UIntToBits_NUM_BITS_64(
	input clk,
	input wire[63:0] value,
	output /*mux_wire*/ logic[63:0] bits
);

	assign bits = value;
endmodule

// BitsToUInt #(NUM_BITS: 11)
module BitsToUInt_NUM_BITS_11(
	input clk,
	input wire[10:0] bits,
	output /*mux_wire*/ logic[10:0] value
);

	assign value = bits;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 4294967296, FROM: 1, TO: 4294967296)
module IntNarrow_FROM_I_0_TO_I_4294967296_FROM_1_TO_4294967296(
	input clk,
	input wire[31:0] in,
	output /*mux_wire*/ logic[31:0] out
);

	assign out = in;
endmodule

// BitsToUInt #(NUM_BITS: 32)
module BitsToUInt_NUM_BITS_32(
	input clk,
	input wire[31:0] bits,
	output /*mux_wire*/ logic[31:0] value
);

	assign value = bits;
endmodule

// axi_memory_writer_tie_off #(AXI_WIDTH: 32)
module axi_memory_writer_tie_off_AXI_WIDTH_32(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic awvalid,
	input wire awready,
	output /*mux_wire*/ logic[63:0] awaddr,
	output /*mux_wire*/ logic[7:0] awlen,
	output /*mux_wire*/ logic[2:0] awsize,
	output /*mux_wire*/ logic[1:0] awburst,
	output /*mux_wire*/ logic[2:0] awprot,
	output /*mux_wire*/ logic[3:0] awcache,
	output /*mux_wire*/ logic[3:0] awqos,
	output /*mux_wire*/ logic awlock,
	output /*mux_wire*/ logic[3:0] awregion,
	output /*mux_wire*/ logic wvalid,
	input wire wready,
	output /*mux_wire*/ logic[31:0] wdata,
	output /*mux_wire*/ logic[3:0] wstrb,
	output /*mux_wire*/ logic wlast,
	input wire bvalid,
	input wire[1:0] bresp,
	output /*mux_wire*/ logic bready
);

/*mux_wire*/ logic _aresetn;
localparam[1:0] _4 = 2'b00;
localparam[2:0] _5 = 3'b000;
localparam[3:0] _6 = 4'b0000;
/*mux_wire*/ logic _Repeat_v;
wire[31:0] _Repeat_result;
/*mux_wire*/ logic _Repeat_2_v;
wire[3:0] _Repeat_2_result;
/*mux_wire*/ logic _awready;
/*mux_wire*/ logic _wready;
/*mux_wire*/ logic _bvalid;
/*mux_wire*/ logic[1:0] _bresp;
Repeat_T_type_bool_SIZE_32 Repeat(
	.clk(aclk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
Repeat_T_type_bool_SIZE_4 Repeat_2(
	.clk(aclk),
	.v(_Repeat_2_v),
	.result(_Repeat_2_result)
);
always_comb begin // combinatorial _aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_aresetn = 1'bx;
	_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_aresetn = _aresetn;
end
always_comb begin // combinatorial awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awvalid = 1'bx;
	awvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awvalid = awvalid;
end
always_comb begin // combinatorial awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awaddr = 64'dx;
	awaddr = 1'd0;
end
always_comb begin // combinatorial awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlen = 8'dx;
	awlen = 1'd0;
end
always_comb begin // combinatorial awsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awsize = 3'dx;
	awsize = 2'd2;
end
always_comb begin // combinatorial awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awburst = 2'bxx;
	awburst = _4;
end
always_comb begin // combinatorial awprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awprot = 3'bxxx;
	awprot = _5;
end
always_comb begin // combinatorial awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awcache = 4'bxxxx;
	awcache = _6;
end
always_comb begin // combinatorial awqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awqos = 4'dx;
	awqos = 1'd0;
end
always_comb begin // combinatorial awlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlock = 1'bx;
	awlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awlock = awlock;
end
always_comb begin // combinatorial awregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awregion = 4'dx;
	awregion = 1'd0;
end
always_comb begin // combinatorial wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wvalid = 1'bx;
	wvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wvalid = wvalid;
end
always_comb begin // combinatorial wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	wdata = _Repeat_result;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	_Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
always_comb begin // combinatorial wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wstrb = 4'bxxxx;
	wstrb = _Repeat_2_result;
end
always_comb begin // combinatorial _Repeat_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_2_v = 1'bx;
	_Repeat_2_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_2_v = _Repeat_2_v;
end
always_comb begin // combinatorial wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wlast = 1'bx;
	wlast = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wlast = wlast;
end
always_comb begin // combinatorial bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	bready = 1'bx;
	bready = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	bready = bready;
end
always_comb begin // combinatorial _awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_awready = 1'bx;
	_awready = awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_awready = _awready;
end
always_comb begin // combinatorial _wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_wready = 1'bx;
	_wready = wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_wready = _wready;
end
always_comb begin // combinatorial _bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_bvalid = 1'bx;
	_bvalid = bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_bvalid = _bvalid;
end
always_comb begin // combinatorial _bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_bresp = 2'bxx;
	_bresp = bresp;
end
endmodule

// axi_realigning_burst_reader #(T: type bool #()[32][1], AXI_WIDTH: 32, ADDR_ALIGN: 4, COUNT_TO: 4294967296, ATO: 18446744073709551616)
module axi_realigning_burst_reader_T_type_bool_32_1_AXI_WIDTH_32_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic arvalid,
	input wire arready,
	output /*mux_wire*/ logic[63:0] araddr,
	output /*mux_wire*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[31:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[31:0] count,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic value_valid,
	output /*mux_wire*/ logic[31:0] value[0:0],
	output /*mux_wire*/ logic last
);

/*mux_wire*/ logic _parent_aresetn;
wire _parent_arvalid;
wire[63:0] _parent_araddr;
wire[7:0] _parent_arlen;
wire[2:0] _parent_arsize;
wire[1:0] _parent_arburst;
wire[2:0] _parent_arprot;
wire[3:0] _parent_arcache;
wire[3:0] _parent_arqos;
wire _parent_arlock;
wire[3:0] _parent_arregion;
wire _parent_rready;
/*mux_wire*/ logic _parent_arready;
/*mux_wire*/ logic _parent_rvalid;
/*mux_wire*/ logic[31:0] _parent_rdata;
/*mux_wire*/ logic[1:0] _parent_rresp;
/*mux_wire*/ logic _parent_rlast;
/*mux_wire*/ logic[10:0] _parent_max_in_flight;
wire _parent_may_request_new_burst;
wire[31:0] _22;
assign _22 = count * 1'd1;
/*mux_wire*/ logic _parent_request_new_burst;
/*mux_wire*/ logic[63:0] _parent_start_addr;
/*mux_wire*/ logic[31:0] _parent_count;
/*mux_wire*/ logic _parent_is_ready_to_receive_lots_of_data;
// (zero sized) stored_elements
// (zero sized) cur_element_store_align
wire _parent_element_packet_valid;
wire[31:0] _parent_elements[0:0];
// (zero sized) _parent_chunk_offset
wire[0:0] _parent_chunk_length;
wire _parent_last;
/*mux_wire*/ logic[31:0] elements[0:0];
// (zero sized) chunk_offset
/*mux_wire*/ logic[0:0] chunk_length;
/*mux_wire*/ logic last_2;
/*mux_wire*/ logic[31:0] elements_extended[0:0];
/*mux_wire*/ logic[31:0] rotated_elements[0:0];
// (zero sized) _31
// (zero sized) _32
/*mux_wire*/ logic[31:0] _RotateRight_data[0:0];
// (zero sized) _RotateRight_offset
wire[31:0] _RotateRight_rotated_data[0:0];
/*mux_wire*/ logic[0:0] rotated_strobe;
// (zero sized) _MakeStrobe_chunk_offset
/*mux_wire*/ logic[0:0] _MakeStrobe_chunk_length;
wire[0:0] _MakeStrobe_strobe;
/*mux_wire*/ logic[0:0] end_of_element;
wire[0:0] _37;
assign _37 = 1'd0 + chunk_length;
wire _39;
assign _39 = end_of_element >= 1'd1;
/*mux_wire*/ logic[31:0] resulting_value_bits;
wire[31:0] _40 = rotated_elements[0];
/*mux_wire*/ logic[31:0] _FromBits_bits;
wire[31:0] _FromBits_value[0:0];
// (zero sized) _45
wire _47;
assign _47 = !aresetn;
axi_array_burst_reader_AXI_WIDTH_32_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616 parent(
	.aclk(aclk),
	.aresetn(_parent_aresetn),
	.arvalid(_parent_arvalid),
	.arready(_parent_arready),
	.araddr(_parent_araddr),
	.arlen(_parent_arlen),
	.arsize(_parent_arsize),
	.arburst(_parent_arburst),
	.arprot(_parent_arprot),
	.arcache(_parent_arcache),
	.arqos(_parent_arqos),
	.arlock(_parent_arlock),
	.arregion(_parent_arregion),
	.rvalid(_parent_rvalid),
	.rready(_parent_rready),
	.rdata(_parent_rdata),
	.rresp(_parent_rresp),
	.rlast(_parent_rlast),
	.is_ready_to_receive_lots_of_data(_parent_is_ready_to_receive_lots_of_data),
	.element_packet_valid(_parent_element_packet_valid),
	.elements(_parent_elements),
	// (zero sized port) .chunk_offset(_parent_chunk_offset)
	.chunk_length(_parent_chunk_length),
	.last(_parent_last),
	.max_in_flight(_parent_max_in_flight),
	.may_request_new_burst(_parent_may_request_new_burst),
	.request_new_burst(_parent_request_new_burst),
	.start_addr(_parent_start_addr),
	.count(_parent_count)
);
RotateRight_T_type_bool_32_ARRAY_LEN_1 RotateRight(
	.clk(aclk),
	.data(_RotateRight_data),
	// (zero sized port) .offset(_RotateRight_offset)
	.rotated_data(_RotateRight_rotated_data)
);
MakeStrobe_STROBE_WIDTH_1 MakeStrobe(
	.clk(aclk),
	// (zero sized port) .chunk_offset(_MakeStrobe_chunk_offset)
	.chunk_length(_MakeStrobe_chunk_length),
	.strobe(_MakeStrobe_strobe)
);
FromBits_T_type_bool_32_1 FromBits(
	.clk(aclk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial _parent_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_aresetn = 1'bx;
	_parent_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_aresetn = _parent_aresetn;
end
always_comb begin // combinatorial arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arvalid = 1'bx;
	arvalid = _parent_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arvalid = arvalid;
end
always_comb begin // combinatorial araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	araddr = 64'dx;
	araddr = _parent_araddr;
end
always_comb begin // combinatorial arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlen = 8'dx;
	arlen = _parent_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = _parent_arsize;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _parent_arburst;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _parent_arprot;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _parent_arcache;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = _parent_arqos;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = _parent_arlock;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = _parent_arregion;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = _parent_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _parent_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_arready = 1'bx;
	_parent_arready = arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_arready = _parent_arready;
end
always_comb begin // combinatorial _parent_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rvalid = 1'bx;
	_parent_rvalid = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rvalid = _parent_rvalid;
end
always_comb begin // combinatorial _parent_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_parent_rdata = rdata;
end
always_comb begin // combinatorial _parent_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rresp = 2'bxx;
	_parent_rresp = rresp;
end
always_comb begin // combinatorial _parent_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rlast = 1'bx;
	_parent_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rlast = _parent_rlast;
end
always_comb begin // combinatorial _parent_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_max_in_flight = 11'dx;
	_parent_max_in_flight = max_in_flight;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _parent_may_request_new_burst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial _parent_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_request_new_burst = 1'bx;
	_parent_request_new_burst = 1'b0;
	if(request_new_burst) _parent_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_request_new_burst = _parent_request_new_burst;
end
always_comb begin // combinatorial _parent_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_start_addr = 64'dx;
	if(request_new_burst) _parent_start_addr = start_addr;
end
always_comb begin // combinatorial _parent_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_count = 32'dx;
	if(request_new_burst) _parent_count = _22;
end
always_comb begin // combinatorial _parent_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_is_ready_to_receive_lots_of_data = 1'bx;
	_parent_is_ready_to_receive_lots_of_data = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_is_ready_to_receive_lots_of_data = _parent_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value_valid = 1'bx;
	value_valid = 1'b0;
	if(_parent_element_packet_valid) if(_39) value_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	value_valid = value_valid;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) value[_v0] = _FromBits_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_parent_element_packet_valid) if(_39) last = last_2;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements[_v0] = _parent_elements[_v0];
end
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 1'dx;
	if(_parent_element_packet_valid) chunk_length = _parent_chunk_length;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunk_length = chunk_length;
end
always_comb begin // combinatorial last_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last_2 = 1'bx;
	if(_parent_element_packet_valid) last_2 = _parent_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last_2 = last_2;
end
always_comb begin // combinatorial elements_extended
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_extended = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements_extended[_v0] = elements[_v0];
end
end
always_comb begin // combinatorial rotated_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) rotated_elements[_v0] = _RotateRight_rotated_data[_v0];
end
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) _RotateRight_data[_v0] = elements_extended[_v0];
end
end
always_comb begin // combinatorial rotated_strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_strobe = 1'bx;
	if(_parent_element_packet_valid) rotated_strobe = _MakeStrobe_strobe;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rotated_strobe = rotated_strobe;
end
always_comb begin // combinatorial _MakeStrobe_chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_length = 1'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_length = chunk_length;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_MakeStrobe_chunk_length = _MakeStrobe_chunk_length;
end
always_comb begin // combinatorial end_of_element
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	end_of_element = 1'dx;
	if(_parent_element_packet_valid) end_of_element = _37;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	end_of_element = end_of_element;
end
always_comb begin // combinatorial resulting_value_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	resulting_value_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) resulting_value_bits[_v0] = _40[_v0];
end
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_parent_element_packet_valid) if(_39) _FromBits_bits = resulting_value_bits;
end
endmodule

// FromBits #(T: type bool #()[32][1])
module FromBits_T_type_bool_32_1(
	input clk,
	input wire[31:0] bits,
	output /*mux_wire*/ logic[31:0] value[0:0]
);

genvar _g0;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign value[_g0] = bits[(_g0) * 32 +: 32];
end
endgenerate
endmodule

// RotateRight #(T: type bool #()[32], ARRAY_LEN: 1)
module RotateRight_T_type_bool_32_ARRAY_LEN_1(
	input clk,
	input wire[31:0] data[0:0],
	// (zero sized) input offset
	output /*mux_wire*/ logic[31:0] rotated_data[0:0]
);

genvar _g0;
// (zero sized) offset_bits
// (zero sized) _UIntToBits_value
// (zero sized) _UIntToBits_bits
/*mux_wire*/ logic[31:0] rotate_stages[0:0][0:0];
wire[31:0] _3[0:0];
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _3[_g0] = rotate_stages[0][_g0];
end
endgenerate
UIntToBits_NUM_BITS_0 UIntToBits(
	.clk(clk)
	// (zero sized port) .value(_UIntToBits_value)
	// (zero sized port) .bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
rotated_data[_v0] = _3[_v0];
end
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{'{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
rotate_stages[0][_v0] = data[_v0];
end
end
endmodule

// axi_array_burst_reader #(AXI_WIDTH: 32, ADDR_ALIGN: 4, COUNT_TO: 4294967296, ATO: 18446744073709551616)
module axi_array_burst_reader_AXI_WIDTH_32_ADDR_ALIGN_4_COUNT_TO_4294967296_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*state*/ logic arvalid,
	input wire arready,
	output /*state*/ logic[63:0] araddr,
	output /*state*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[31:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic element_packet_valid,
	output /*mux_wire*/ logic[31:0] elements[0:0],
	// (zero sized) output chunk_offset
	output /*mux_wire*/ logic[0:0] chunk_length,
	output /*mux_wire*/ logic last,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[31:0] count
);

/*latency*/ logic _arvalid_D1; always_ff @(posedge aclk) begin _arvalid_D1 <= arvalid; end
/*latency*/ logic _request_new_burst_D1; always_ff @(posedge aclk) begin _request_new_burst_D1 <= request_new_burst; end
genvar _g0;
localparam[1:0] _1 = 2'b01;
localparam[2:0] _2 = 3'b000;
localparam[3:0] _3 = 4'b0010;
/*mux_wire*/ logic[1:0] _rresp;
/*mux_wire*/ logic _rlast;
/*state*/ logic[11:0] num_in_flight;
/*state*/ logic last_burst_in_flight;
/*mux_wire*/ logic[63:0] next_araddr;
/*latency*/ logic[63:0] _next_araddr_D0; always_ff @(posedge aclk) begin _next_araddr_D0 <= next_araddr; end
wire[61:0] _cur_start_chunk_addr_old;
/*mux_wire*/ logic[61:0] _BitwiseIntConcat_upper;
/*mux_wire*/ logic[1:0] _BitwiseIntConcat_lower;
wire[63:0] _BitwiseIntConcat_v;
/*mux_wire*/ logic[7:0] next_arlen;
/*mux_wire*/ logic next_last_burst_in_flight;
/*latency*/ logic _next_last_burst_in_flight_D0; always_ff @(posedge aclk) begin _next_last_burst_in_flight_D0 <= next_last_burst_in_flight; end
/*mux_wire*/ logic[53:0] cur_burst_addr;
/*mux_wire*/ logic[7:0] cur_align;
/*mux_wire*/ logic[61:0] _BitwiseIntSplit_v;
wire[53:0] _BitwiseIntSplit_upper;
wire[7:0] _BitwiseIntSplit_lower;
/*mux_wire*/ logic chunks_are_left;
/*latency*/ logic _chunks_are_left_D0; always_ff @(posedge aclk) begin _chunks_are_left_D0 <= chunks_are_left; end
wire[32:0] _num_chunks_left_old;
/*latency*/ logic[32:0] __num_chunks_left_old_N1; always_ff @(posedge aclk) begin __num_chunks_left_old_N1 <= _num_chunks_left_old; end
/*latency*/ logic[32:0] __num_chunks_left_old_D0; always_ff @(posedge aclk) begin __num_chunks_left_old_D0 <= __num_chunks_left_old_N1; end
wire _14;
assign _14 = _num_chunks_left_old > 1'd0;
/*latency*/ logic __14_N1; always_ff @(posedge aclk) begin __14_N1 <= _14; end
/*mux_wire*/ logic[7:0] max_chunks_in_this_burst;
/*latency*/ logic[7:0] _max_chunks_in_this_burst_D0; always_ff @(posedge aclk) begin _max_chunks_in_this_burst_D0 <= max_chunks_in_this_burst; end
wire[7:0] _18;
assign _18 = 8'd255 - cur_align;
wire[8:0] _22;
assign _22 = max_chunks_in_this_burst + 1'd1;
wire _23;
assign _23 = __num_chunks_left_old_N1 <= _22;
/*latency*/ logic __23_D0; always_ff @(posedge aclk) begin __23_D0 <= _23; end
/*mux_wire*/ logic[32:0] _IntNarrow_in;
wire[8:0] _IntNarrow_out;
wire[7:0] _26;
assign _26 = _IntNarrow_out - 1'd1;
/*latency*/ logic[7:0] __26_D0; always_ff @(posedge aclk) begin __26_D0 <= _26; end
/*mux_wire*/ logic may_next_arvalid;
/*latency*/ logic _may_next_arvalid_D1; always_ff @(posedge aclk) begin _may_next_arvalid_D1 <= may_next_arvalid; end
wire _num_chunks_left_may_update;
wire _30;
assign _30 = _chunks_are_left_D0 & _num_chunks_left_may_update;
wire _cur_start_chunk_addr_may_update;
wire _32;
assign _32 = _30 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
wire _34;
assign _34 = _32 & _LatencyOffset_out;
wire signed[11:0] _37;
assign _37 = max_in_flight - 9'd256;
wire _38;
assign _38 = $signed({1'b0, num_in_flight}) <= _37;
wire _39;
assign _39 = _34 & _38;
/*mux_wire*/ logic[54:0] next_burst_addr;
wire[54:0] _45;
assign _45 = cur_burst_addr + 1'd1;
/*latency*/ logic[54:0] __45_D0; always_ff @(posedge aclk) begin __45_D0 <= _45; end
/*latency*/ logic[54:0] __45_D1; always_ff @(posedge aclk) begin __45_D1 <= __45_D0; end
/*mux_wire*/ logic[54:0] _BitwiseIntConcat_2_upper;
/*mux_wire*/ logic[7:0] _BitwiseIntConcat_2_lower;
wire[62:0] _BitwiseIntConcat_2_v;
/*mux_wire*/ logic[62:0] _IntNarrow_2_in;
wire[61:0] _IntNarrow_2_out;
/*mux_wire*/ logic _cur_start_chunk_addr_update;
/*mux_wire*/ logic[61:0] _cur_start_chunk_addr_new;
/*mux_wire*/ logic[32:0] next_num_chunks_left;
wire[8:0] _53;
assign _53 = next_arlen + 1'd1;
wire signed[33:0] _54;
assign _54 = __num_chunks_left_old_D0 - _53;
/*mux_wire*/ logic signed[33:0] _IntNarrow_3_in;
wire[32:0] _IntNarrow_3_out;
/*mux_wire*/ logic _num_chunks_left_update;
/*mux_wire*/ logic[32:0] _num_chunks_left_new;
/*mux_wire*/ logic _BoolToInt_i;
wire[0:0] _BoolToInt_o;
wire signed[12:0] _64;
assign _64 = num_in_flight - _BoolToInt_o;
wire _66;
assign _66 = !arvalid;
wire _68;
assign _68 = _66 & may_next_arvalid;
wire[8:0] _71;
assign _71 = next_arlen + 1'd1;
/*mux_wire*/ logic _Ternary_cond;
/*mux_wire*/ logic[8:0] _Ternary_a;
/*mux_wire*/ logic[8:0] _Ternary_b;
wire[8:0] _Ternary_o;
wire signed[12:0] _73;
assign _73 = _64 + $signed({1'b0, _Ternary_o});
/*mux_wire*/ logic signed[12:0] _IntNarrow_4_in;
wire[11:0] _IntNarrow_4_out;
/*state*/ logic[0:0] final_chunk_align;
// (zero sized) cur_chunk_align
/*mux_wire*/ logic[31:0] elements_2[0:0];
wire[31:0] _75;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _75[_g0] = rdata[_g0];
end
endgenerate
/*mux_wire*/ logic[0:0] num_chunk_elements;
/*mux_wire*/ logic is_last;
wire _78;
assign _78 = num_in_flight == 1'd1;
wire _80;
assign _80 = _78 & last_burst_in_flight;
wire[0:0] _84;
assign _84 = final_chunk_align - 1'd0;
/*mux_wire*/ logic[0:0] _IntNarrow_5_in;
wire[0:0] _IntNarrow_5_out;
wire[0:0] _86;
assign _86 = 1'd1 - 1'd0;
wire _94;
assign _94 = !chunks_are_left;
/*latency*/ logic __94_D0; always_ff @(posedge aclk) begin __94_D0 <= _94; end
wire _96;
assign _96 = __94_D0 & _num_chunks_left_may_update;
wire _98;
assign _98 = _96 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic[61:0] chunk_addr;
/*latency*/ logic[61:0] _chunk_addr_D1; always_ff @(posedge aclk) begin _chunk_addr_D1 <= chunk_addr; end
// (zero sized) element_in_chunk_align
wire[61:0] _100;
assign _100 = start_addr / 3'd4;
/*mux_wire*/ logic[61:0] _BitwiseIntSplit_2_v;
wire[61:0] _BitwiseIntSplit_2_upper;
// (zero sized) _BitwiseIntSplit_2_lower
/*mux_wire*/ logic[31:0] chunk_count_bits;
// (zero sized) final_alignment
wire[31:0] _103;
assign _103 = count + 1'd0;
/*mux_wire*/ logic[31:0] _BitwiseIntSplit_3_v;
wire[31:0] _BitwiseIntSplit_3_upper;
// (zero sized) _BitwiseIntSplit_3_lower
/*mux_wire*/ logic[32:0] num_chunks;
/*mux_wire*/ logic is_no_chunks;
wire _106;
assign _106 = chunk_count_bits == 1'd0;
wire _112;
assign _112 = 1'd0 != 1'd0;
/*mux_wire*/ logic _BoolToInt_2_i;
wire[0:0] _BoolToInt_2_o;
wire[32:0] _113;
assign _113 = chunk_count_bits + _BoolToInt_2_o;
wire _119;
assign _119 = !is_no_chunks;
wire _122;
assign _122 = 1'd0 == 1'd0;
wire _123;
assign _123 = _119 & _122;
/*mux_wire*/ logic _BoolToInt_3_i;
wire[0:0] _BoolToInt_3_o;
/*mux_wire*/ logic[0:0] _BitwiseIntConcat_3_upper;
// (zero sized) _BitwiseIntConcat_3_lower
wire[0:0] _BitwiseIntConcat_3_v;
wire _127;
assign _127 = !aresetn;
/*mux_wire*/ logic _cur_start_chunk_addr_rst;
wire _129;
assign _129 = !aresetn;
/*mux_wire*/ logic _num_chunks_left_rst;
wire _131;
assign _131 = !aresetn;
SlowState_T_type_int_FROM_0_TO_4611686018427387904_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1 cur_start_chunk_addr(
	.clk(aclk),
	.rst(_cur_start_chunk_addr_rst),
	.old(_cur_start_chunk_addr_old),
	.may_update(_cur_start_chunk_addr_may_update),
	.update(_cur_start_chunk_addr_update),
	.new_1(_cur_start_chunk_addr_new)
);
SlowState_T_type_int_FROM_0_TO_4294967299_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0 num_chunks_left(
	.clk(aclk),
	.rst(_num_chunks_left_rst),
	.old(_num_chunks_left_old),
	.may_update(_num_chunks_left_may_update),
	.update(_num_chunks_left_update),
	.new_1(_num_chunks_left_new)
);
BitwiseIntConcat_UPPER_TO_4611686018427387904_LOWER_BITS_2 BitwiseIntConcat(
	.clk(aclk),
	.upper(_BitwiseIntConcat_upper),
	.lower(_BitwiseIntConcat_lower),
	.v(_BitwiseIntConcat_v)
);
BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_8 BitwiseIntSplit(
	.clk(aclk),
	.v(_BitwiseIntSplit_v),
	.upper(_BitwiseIntSplit_upper),
	.lower(_BitwiseIntSplit_lower)
);
IntNarrow_FROM_I_0_TO_I_4294967299_FROM_1_TO_257 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
LatencyOffset_T_type_bool_OFFSET_384 LatencyOffset(
	.clk(aclk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
BitwiseIntConcat_UPPER_TO_18014398509481985_LOWER_BITS_8 BitwiseIntConcat_2(
	.clk(aclk),
	.upper(_BitwiseIntConcat_2_upper),
	.lower(_BitwiseIntConcat_2_lower),
	.v(_BitwiseIntConcat_2_v)
);
IntNarrow_FROM_I_0_TO_I_4611686018427388160_FROM_0_TO_4611686018427387904 IntNarrow_2(
	.clk(aclk),
	.in(_IntNarrow_2_in),
	.out(_IntNarrow_2_out)
);
IntNarrow_FROM_I_256_TO_I_4294967298_FROM_0_TO_4294967299 IntNarrow_3(
	.clk(aclk),
	.in(_IntNarrow_3_in),
	.out(_IntNarrow_3_out)
);
BoolToInt BoolToInt(
	.clk(aclk),
	.i(_BoolToInt_i),
	.o(_BoolToInt_o)
);
Ternary_T_type_int_FROM_0_TO_257 Ternary(
	.clk(aclk),
	.cond(_Ternary_cond),
	.a(_Ternary_a),
	.b(_Ternary_b),
	.o(_Ternary_o)
);
IntNarrow_FROM_I_1_TO_I_3640_FROM_0_TO_3384 IntNarrow_4(
	.clk(aclk),
	.in(_IntNarrow_4_in),
	.out(_IntNarrow_4_out)
);
IntNarrow_FROM_I_0_TO_I_2_FROM_0_TO_2 IntNarrow_5(
	.clk(aclk),
	.in(_IntNarrow_5_in),
	.out(_IntNarrow_5_out)
);
BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_0 BitwiseIntSplit_2(
	.clk(aclk),
	.v(_BitwiseIntSplit_2_v),
	.upper(_BitwiseIntSplit_2_upper)
	// (zero sized port) .lower(_BitwiseIntSplit_2_lower)
);
BitwiseIntSplit_TO_4294967296_LOWER_BITS_0 BitwiseIntSplit_3(
	.clk(aclk),
	.v(_BitwiseIntSplit_3_v),
	.upper(_BitwiseIntSplit_3_upper)
	// (zero sized port) .lower(_BitwiseIntSplit_3_lower)
);
BoolToInt BoolToInt_2(
	.clk(aclk),
	.i(_BoolToInt_2_i),
	.o(_BoolToInt_2_o)
);
BoolToInt BoolToInt_3(
	.clk(aclk),
	.i(_BoolToInt_3_i),
	.o(_BoolToInt_3_o)
);
BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_0 BitwiseIntConcat_3(
	.clk(aclk),
	.upper(_BitwiseIntConcat_3_upper),
	// (zero sized port) .lower(_BitwiseIntConcat_3_lower)
	.v(_BitwiseIntConcat_3_v)
);
always_ff @(posedge aclk) begin // state arvalid
	if(arvalid) if(arready) arvalid <= 1'b0;
	if(!arvalid) if(may_next_arvalid) arvalid <= 1'b1;
	if(_131) arvalid <= 1'b0;
end
always_ff @(posedge aclk) begin // state araddr
	if(!arvalid) if(may_next_arvalid) araddr <= _next_araddr_D0;
end
always_ff @(posedge aclk) begin // state arlen
	if(!arvalid) if(may_next_arvalid) arlen <= next_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = 2'd2;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _1;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _2;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _3;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = 1'd0;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = 1'd0;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rresp = 2'bxx;
	_rresp = rresp;
end
always_comb begin // combinatorial _rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rlast = 1'bx;
	_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_rlast = _rlast;
end
always_comb begin // combinatorial element_packet_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_packet_valid = 1'bx;
	element_packet_valid = 1'b0;
	if(rvalid) element_packet_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	element_packet_valid = element_packet_valid;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(rvalid) elements[_v0] = elements_2[_v0];
end
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 1'dx;
	if(rvalid) chunk_length = num_chunk_elements;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunk_length = chunk_length;
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(rvalid) last = is_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state num_in_flight
	num_in_flight <= _IntNarrow_4_out;
	if(_131) num_in_flight <= 1'd0;
end
always_ff @(posedge aclk) begin // state last_burst_in_flight
	if(!arvalid) if(may_next_arvalid) last_burst_in_flight <= _next_last_burst_in_flight_D0;
end
always_comb begin // combinatorial next_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_araddr = 64'dx;
	next_araddr = _BitwiseIntConcat_v;
end
always_comb begin // combinatorial _BitwiseIntConcat_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_upper = 62'dx;
	_BitwiseIntConcat_upper = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial _BitwiseIntConcat_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_lower = 2'dx;
	_BitwiseIntConcat_lower = 1'd0;
end
always_comb begin // combinatorial next_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_arlen = 8'dx;
	if(_chunks_are_left_D0) if(__23_D0) next_arlen = __26_D0;
	if(_chunks_are_left_D0) if(!__23_D0) next_arlen = _max_chunks_in_this_burst_D0;
end
always_comb begin // combinatorial next_last_burst_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_last_burst_in_flight = 1'bx;
	next_last_burst_in_flight = 1'b0;
	if(chunks_are_left) if(_23) next_last_burst_in_flight = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	next_last_burst_in_flight = next_last_burst_in_flight;
end
always_comb begin // combinatorial cur_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_burst_addr = 54'dx;
	cur_burst_addr = _BitwiseIntSplit_upper;
end
always_comb begin // combinatorial cur_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_align = 8'dx;
	cur_align = _BitwiseIntSplit_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_v = 62'dx;
	_BitwiseIntSplit_v = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial chunks_are_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunks_are_left = 1'bx;
	chunks_are_left = __14_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunks_are_left = chunks_are_left;
end
always_comb begin // combinatorial max_chunks_in_this_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	max_chunks_in_this_burst = 8'dx;
	if(chunks_are_left) max_chunks_in_this_burst = _18;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 33'dx;
	if(chunks_are_left) if(_23) _IntNarrow_in = __num_chunks_left_old_N1;
end
always_comb begin // combinatorial may_next_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_next_arvalid = 1'bx;
	may_next_arvalid = _39;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_next_arvalid = may_next_arvalid;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial next_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_burst_addr = 55'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) next_burst_addr = __45_D1;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_upper = 55'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_upper = next_burst_addr;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_lower = 8'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_lower = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_2_in = 63'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _IntNarrow_2_in = _BitwiseIntConcat_2_v;
end
always_comb begin // combinatorial _cur_start_chunk_addr_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_update = 1'bx;
	_cur_start_chunk_addr_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _cur_start_chunk_addr_update = 1'b1;
	if(request_new_burst) _cur_start_chunk_addr_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_update = _cur_start_chunk_addr_update;
end
always_comb begin // combinatorial _cur_start_chunk_addr_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_new = 62'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _cur_start_chunk_addr_new = _IntNarrow_2_out;
	if(_request_new_burst_D1) _cur_start_chunk_addr_new = _chunk_addr_D1;
end
always_comb begin // combinatorial next_num_chunks_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_num_chunks_left = 33'dx;
	if(!arvalid) if(may_next_arvalid) next_num_chunks_left = _IntNarrow_3_out;
end
always_comb begin // combinatorial _IntNarrow_3_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_3_in = 34'sdx;
	if(!arvalid) if(may_next_arvalid) _IntNarrow_3_in = _54;
end
always_comb begin // combinatorial _num_chunks_left_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_update = 1'bx;
	_num_chunks_left_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_update = 1'b1;
	if(request_new_burst) _num_chunks_left_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_update = _num_chunks_left_update;
end
always_comb begin // combinatorial _num_chunks_left_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_new = 33'dx;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_new = next_num_chunks_left;
	if(request_new_burst) _num_chunks_left_new = num_chunks;
end
always_comb begin // combinatorial _BoolToInt_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_i = 1'bx;
	_BoolToInt_i = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_i = _BoolToInt_i;
end
always_comb begin // combinatorial _Ternary_cond
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_cond = 1'bx;
	_Ternary_cond = _68;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Ternary_cond = _Ternary_cond;
end
always_comb begin // combinatorial _Ternary_a
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_a = 9'dx;
	_Ternary_a = _71;
end
always_comb begin // combinatorial _Ternary_b
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_b = 9'dx;
	_Ternary_b = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_4_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_4_in = 13'sdx;
	_IntNarrow_4_in = _73;
end
always_ff @(posedge aclk) begin // state final_chunk_align
	if(request_new_burst) final_chunk_align <= _BitwiseIntConcat_3_v;
end
always_comb begin // combinatorial elements_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_2 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	if(rvalid) elements_2[0] = _75;
end
always_comb begin // combinatorial num_chunk_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunk_elements = 1'dx;
	if(rvalid) if(is_last) num_chunk_elements = _IntNarrow_5_out;
	if(rvalid) if(!is_last) num_chunk_elements = _86;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	num_chunk_elements = num_chunk_elements;
end
always_comb begin // combinatorial is_last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_last = 1'bx;
	if(rvalid) is_last = _80;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_last = is_last;
end
always_comb begin // combinatorial _IntNarrow_5_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_5_in = 1'dx;
	if(rvalid) if(is_last) _IntNarrow_5_in = _84;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_IntNarrow_5_in = _IntNarrow_5_in;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _98;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial chunk_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_addr = 62'dx;
	if(request_new_burst) chunk_addr = _BitwiseIntSplit_2_upper;
end
always_comb begin // combinatorial _BitwiseIntSplit_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_2_v = 62'dx;
	if(request_new_burst) _BitwiseIntSplit_2_v = _100;
end
always_comb begin // combinatorial chunk_count_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_count_bits = 32'dx;
	if(request_new_burst) chunk_count_bits = _BitwiseIntSplit_3_upper;
end
always_comb begin // combinatorial _BitwiseIntSplit_3_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_3_v = 32'dx;
	if(request_new_burst) _BitwiseIntSplit_3_v = _103;
end
always_comb begin // combinatorial num_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunks = 33'dx;
	if(request_new_burst) if(is_no_chunks) num_chunks = 1'd1;
	if(request_new_burst) if(!is_no_chunks) num_chunks = _113;
end
always_comb begin // combinatorial is_no_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_no_chunks = 1'bx;
	if(request_new_burst) is_no_chunks = _106;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_no_chunks = is_no_chunks;
end
always_comb begin // combinatorial _BoolToInt_2_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_2_i = 1'bx;
	if(request_new_burst) if(!is_no_chunks) _BoolToInt_2_i = _112;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_2_i = _BoolToInt_2_i;
end
always_comb begin // combinatorial _BoolToInt_3_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_3_i = 1'bx;
	if(request_new_burst) _BoolToInt_3_i = _123;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_3_i = _BoolToInt_3_i;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_upper = 1'dx;
	if(request_new_burst) _BitwiseIntConcat_3_upper = _BoolToInt_3_o;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BitwiseIntConcat_3_upper = _BitwiseIntConcat_3_upper;
end
always_comb begin // combinatorial _cur_start_chunk_addr_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_rst = 1'bx;
	_cur_start_chunk_addr_rst = _127;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_rst = _cur_start_chunk_addr_rst;
end
always_comb begin // combinatorial _num_chunks_left_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_rst = 1'bx;
	_num_chunks_left_rst = _129;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_rst = _num_chunks_left_rst;
end
endmodule

// BitwiseIntSplit #(TO: 4294967296, LOWER_BITS: 0)
module BitwiseIntSplit_TO_4294967296_LOWER_BITS_0(
	input clk,
	input wire[31:0] v,
	output /*mux_wire*/ logic[31:0] upper
	// (zero sized) output lower
);

genvar _g0;
/*mux_wire*/ logic[31:0] v_bits;
/*mux_wire*/ logic[31:0] _UIntToBits_value;
wire[31:0] _UIntToBits_bits;
// (zero sized) _2
// (zero sized) _BitsToUInt_bits
// (zero sized) _BitsToUInt_value
wire[31:0] _3;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[31:0] _FromBits_bits;
wire[31:0] _FromBits_value;
UIntToBits_NUM_BITS_32 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_0 BitsToUInt(
	.clk(clk)
	// (zero sized port) .bits(_BitsToUInt_bits)
	// (zero sized port) .value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_4294967296 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 32'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 32'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 4294967296))
module FromBits_T_type_int_FROM_0_TO_4294967296(
	input clk,
	input wire[31:0] bits,
	output /*mux_wire*/ logic[31:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 32)
module UIntToBits_NUM_BITS_32(
	input clk,
	input wire[31:0] value,
	output /*mux_wire*/ logic[31:0] bits
);

	assign bits = value;
endmodule

// BitwiseIntSplit #(TO: 4611686018427387904, LOWER_BITS: 0)
module BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_0(
	input clk,
	input wire[61:0] v,
	output /*mux_wire*/ logic[61:0] upper
	// (zero sized) output lower
);

genvar _g0;
/*mux_wire*/ logic[61:0] v_bits;
/*mux_wire*/ logic[61:0] _UIntToBits_value;
wire[61:0] _UIntToBits_bits;
// (zero sized) _2
// (zero sized) _BitsToUInt_bits
// (zero sized) _BitsToUInt_value
wire[61:0] _3;
generate
for(_g0 = 0; _g0 < 62; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[61:0] _FromBits_bits;
wire[61:0] _FromBits_value;
UIntToBits_NUM_BITS_62 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_0 BitsToUInt(
	.clk(clk)
	// (zero sized port) .bits(_BitsToUInt_bits)
	// (zero sized port) .value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_4611686018427387904 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 62'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 62'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 62'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 62'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 4611686018427387904))
module FromBits_T_type_int_FROM_0_TO_4611686018427387904(
	input clk,
	input wire[61:0] bits,
	output /*mux_wire*/ logic[61:0] value
);

assign value = bits;
endmodule

// IntNarrow #(FROM_I: -256, TO_I: 4294967298, FROM: 0, TO: 4294967299)
module IntNarrow_FROM_I_256_TO_I_4294967298_FROM_0_TO_4294967299(
	input clk,
	input wire signed[33:0] in,
	output /*mux_wire*/ logic[32:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 4611686018427388160, FROM: 0, TO: 4611686018427387904)
module IntNarrow_FROM_I_0_TO_I_4611686018427388160_FROM_0_TO_4611686018427387904(
	input clk,
	input wire[62:0] in,
	output /*mux_wire*/ logic[61:0] out
);

	assign out = in;
endmodule

// BitwiseIntConcat #(UPPER_TO: 18014398509481985, LOWER_BITS: 8)
module BitwiseIntConcat_UPPER_TO_18014398509481985_LOWER_BITS_8(
	input clk,
	input wire[54:0] upper,
	input wire[7:0] lower,
	output /*mux_wire*/ logic[62:0] v
);

/*mux_wire*/ logic[62:0] v_bits;
/*mux_wire*/ logic[7:0] _UIntToBits_value;
wire[7:0] _UIntToBits_bits;
/*mux_wire*/ logic[54:0] _UIntToBits_2_value;
wire[54:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[62:0] _FromBits_bits;
wire[62:0] _FromBits_value;
UIntToBits_NUM_BITS_8 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_55 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_4611686018427388160 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 63'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 63'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 55; _v0 = _v0 + 1) begin
v_bits[8 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 8'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 55'dx;
	_UIntToBits_2_value = upper;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 63'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 4611686018427388160))
module FromBits_T_type_int_FROM_0_TO_4611686018427388160(
	input clk,
	input wire[62:0] bits,
	output /*mux_wire*/ logic[62:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 55)
module UIntToBits_NUM_BITS_55(
	input clk,
	input wire[54:0] value,
	output /*mux_wire*/ logic[54:0] bits
);

	assign bits = value;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 4294967299, FROM: 1, TO: 257)
module IntNarrow_FROM_I_0_TO_I_4294967299_FROM_1_TO_257(
	input clk,
	input wire[32:0] in,
	output /*mux_wire*/ logic[8:0] out
);

	assign out = in;
endmodule

// BitwiseIntSplit #(TO: 4611686018427387904, LOWER_BITS: 8)
module BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_8(
	input clk,
	input wire[61:0] v,
	output /*mux_wire*/ logic[53:0] upper,
	output /*mux_wire*/ logic[7:0] lower
);

genvar _g0;
/*mux_wire*/ logic[61:0] v_bits;
/*mux_wire*/ logic[61:0] _UIntToBits_value;
wire[61:0] _UIntToBits_bits;
wire[7:0] _2;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[7:0] _BitsToUInt_bits;
wire[7:0] _BitsToUInt_value;
wire[53:0] _3;
generate
for(_g0 = 0; _g0 < 54; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[8 + _g0];
end
endgenerate
/*mux_wire*/ logic[53:0] _FromBits_bits;
wire[53:0] _FromBits_value;
UIntToBits_NUM_BITS_62 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_8 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_18014398509481984 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 54'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 8'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 62'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 62'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 8'bxxxxxxxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 54'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 18014398509481984))
module FromBits_T_type_int_FROM_0_TO_18014398509481984(
	input clk,
	input wire[53:0] bits,
	output /*mux_wire*/ logic[53:0] value
);

assign value = bits;
endmodule

// BitwiseIntConcat #(UPPER_TO: 4611686018427387904, LOWER_BITS: 2)
module BitwiseIntConcat_UPPER_TO_4611686018427387904_LOWER_BITS_2(
	input clk,
	input wire[61:0] upper,
	input wire[1:0] lower,
	output /*mux_wire*/ logic[63:0] v
);

/*mux_wire*/ logic[63:0] v_bits;
/*mux_wire*/ logic[1:0] _UIntToBits_value;
wire[1:0] _UIntToBits_bits;
/*mux_wire*/ logic[61:0] _UIntToBits_2_value;
wire[61:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[63:0] _FromBits_bits;
wire[63:0] _FromBits_value;
UIntToBits_NUM_BITS_2 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_62 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_18446744073709551616 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 64'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 62; _v0 = _v0 + 1) begin
v_bits[2 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 2'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 62'dx;
	_UIntToBits_2_value = upper;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// SlowState #(T: type int #(FROM: 0, TO: 4294967299), RESET_TO: 0, OLD_DELAY: 2, NEW_DELAY: 0)
module SlowState_T_type_int_FROM_0_TO_4294967299_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0(
	input clk,
	input wire rst,
	output /*state*/ logic[32:0] old,
	output /*mux_wire*/ logic may_update,
	input wire update,
	input wire[32:0] new_1
);

genvar _g0;
/*mux_wire*/ logic _cross_rst_in;
/*mux_wire*/ logic[32:0] new_s;
/*mux_wire*/ logic update_s;
/*mux_wire*/ logic update_old;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
/*mux_wire*/ logic[32:0] new_old;
/*mux_wire*/ logic[32:0] _LatencyOffset_2_in;
wire[32:0] _LatencyOffset_2_out;
wire _cross_rst_out;
/*latency*/ logic __cross_rst_out_N1; always_ff @(posedge clk) begin __cross_rst_out_N1 <= _cross_rst_out; end
/*latency*/ logic __cross_rst_out_D0; always_ff @(posedge clk) begin __cross_rst_out_D0 <= __cross_rst_out_N1; end
/*state*/ logic[1:0] cooldown;
wire _8 = cooldown[0];
wire _11;
assign _11 = update_s | __cross_rst_out_D0;
/*mux_wire*/ logic _Repeat_v;
wire[1:0] _Repeat_result;
wire[0:0] _12;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _12[_g0] = cooldown[1 + _g0];
end
endgenerate
CrossDomain_T_type_bool cross_rst(
	.in_clk(clk),
	.in(_cross_rst_in),
	.out(_cross_rst_out)
);
LatencyOffset_T_type_bool_OFFSET_2 LatencyOffset(
	.clk(clk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
LatencyOffset_T_type_int_FROM_0_TO_4294967299_OFFSET_2 LatencyOffset_2(
	.clk(clk),
	.in(_LatencyOffset_2_in),
	.out(_LatencyOffset_2_out)
);
Repeat_T_type_bool_SIZE_2 Repeat(
	.clk(clk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
always_comb begin // combinatorial _cross_rst_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_rst_in = 1'bx;
	_cross_rst_in = rst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_rst_in = _cross_rst_in;
end
always_ff @(posedge clk) begin // state old
	if(_cross_rst_out) old <= 33'd0;
	if(!_cross_rst_out) if(update_old) old <= new_old;
end
always_comb begin // combinatorial new_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_s = 33'dx;
	if(update) new_s = new_1;
end
always_comb begin // combinatorial update_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_s = 1'bx;
	if(update) update_s = 1'b1;
	if(!update) update_s = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_s = update_s;
end
always_comb begin // combinatorial update_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_old = 1'bx;
	update_old = _LatencyOffset_out;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_old = update_old;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = update_s;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial new_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_old = 33'dx;
	new_old = _LatencyOffset_2_out;
end
always_comb begin // combinatorial _LatencyOffset_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_2_in = 33'dx;
	_LatencyOffset_2_in = new_s;
end
always_comb begin // combinatorial may_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_update = 1'bx;
	may_update = _8;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_update = may_update;
end
always_ff @(posedge clk) begin // state cooldown
	if(_11) cooldown <= _Repeat_result;
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(!_11) cooldown[_v0] <= _12[_v0];
end
	if(!_11) cooldown[1] <= 1'b1;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	if(_11) _Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
endmodule

// LatencyOffset #(T: type int #(FROM: 0, TO: 4294967299), OFFSET: -2)
module LatencyOffset_T_type_int_FROM_0_TO_4294967299_OFFSET_2(
	input clk,
	input wire[32:0] in,
	output /*mux_wire*/ logic[32:0] out
);

	assign out = in;
endmodule

// SlowState #(T: type int #(FROM: 0, TO: 4611686018427387904), RESET_TO: 0, OLD_DELAY: 1, NEW_DELAY: 1)
module SlowState_T_type_int_FROM_0_TO_4611686018427387904_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1(
	input clk,
	input wire rst,
	output /*state*/ logic[61:0] old,
	output /*mux_wire*/ logic may_update,
	input wire update,
	input wire[61:0] new_1
);

/*latency*/ logic _update_D1; always_ff @(posedge clk) begin _update_D1 <= update; end
genvar _g0;
/*mux_wire*/ logic _cross_rst_in;
/*mux_wire*/ logic[61:0] new_s;
/*mux_wire*/ logic update_s;
/*mux_wire*/ logic update_old;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
/*latency*/ logic __LatencyOffset_out_N1; always_ff @(posedge clk) begin __LatencyOffset_out_N1 <= _LatencyOffset_out; end
/*mux_wire*/ logic[61:0] new_old;
/*mux_wire*/ logic[61:0] _LatencyOffset_2_in;
wire[61:0] _LatencyOffset_2_out;
wire _cross_rst_out;
/*latency*/ logic __cross_rst_out_D0; always_ff @(posedge clk) begin __cross_rst_out_D0 <= _cross_rst_out; end
/*state*/ logic[1:0] cooldown;
wire _8 = cooldown[0];
wire _11;
assign _11 = update_s | __cross_rst_out_D0;
/*mux_wire*/ logic _Repeat_v;
wire[1:0] _Repeat_result;
wire[0:0] _12;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _12[_g0] = cooldown[1 + _g0];
end
endgenerate
CrossDomain_T_type_bool cross_rst(
	.in_clk(clk),
	.in(_cross_rst_in),
	.out(_cross_rst_out)
);
LatencyOffset_T_type_bool_OFFSET_2 LatencyOffset(
	.clk(clk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
LatencyOffset_T_type_int_FROM_0_TO_4611686018427387904_OFFSET_2 LatencyOffset_2(
	.clk(clk),
	.in(_LatencyOffset_2_in),
	.out(_LatencyOffset_2_out)
);
Repeat_T_type_bool_SIZE_2 Repeat(
	.clk(clk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
always_comb begin // combinatorial _cross_rst_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_rst_in = 1'bx;
	_cross_rst_in = rst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_rst_in = _cross_rst_in;
end
always_ff @(posedge clk) begin // state old
	if(_cross_rst_out) old <= 62'd0;
	if(!_cross_rst_out) if(update_old) old <= new_old;
end
always_comb begin // combinatorial new_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_s = 62'dx;
	if(_update_D1) new_s = new_1;
end
always_comb begin // combinatorial update_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_s = 1'bx;
	if(update) update_s = 1'b1;
	if(!update) update_s = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_s = update_s;
end
always_comb begin // combinatorial update_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_old = 1'bx;
	update_old = __LatencyOffset_out_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_old = update_old;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = update_s;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial new_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_old = 62'dx;
	new_old = _LatencyOffset_2_out;
end
always_comb begin // combinatorial _LatencyOffset_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_2_in = 62'dx;
	_LatencyOffset_2_in = new_s;
end
always_comb begin // combinatorial may_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_update = 1'bx;
	may_update = _8;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_update = may_update;
end
always_ff @(posedge clk) begin // state cooldown
	if(_11) cooldown <= _Repeat_result;
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(!_11) cooldown[_v0] <= _12[_v0];
end
	if(!_11) cooldown[1] <= 1'b1;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	if(_11) _Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
endmodule

// LatencyOffset #(T: type int #(FROM: 0, TO: 4611686018427387904), OFFSET: -2)
module LatencyOffset_T_type_int_FROM_0_TO_4611686018427387904_OFFSET_2(
	input clk,
	input wire[61:0] in,
	output /*mux_wire*/ logic[61:0] out
);

	assign out = in;
endmodule

// axi_ctrl_slave #(NUM_INPUT_REGS: 4, NUM_OUTPUT_REGS: 6, ADDR_WIDTH: 12, AXI_WIDTH: 32)
module axi_ctrl_slave_NUM_INPUT_REGS_4_NUM_OUTPUT_REGS_6_ADDR_WIDTH_12_AXI_WIDTH_32(
	input aclk,
	input wire aresetn,
	input wire[11:0] awaddr,
	input wire awvalid,
	output /*mux_wire*/ logic awready,
	input wire[31:0] wdata,
	input wire[3:0] wstrb,
	input wire wvalid,
	output /*mux_wire*/ logic wready,
	output /*mux_wire*/ logic[1:0] bresp,
	output /*mux_wire*/ logic bvalid,
	input wire bready,
	input wire[11:0] araddr,
	input wire arvalid,
	output /*mux_wire*/ logic arready,
	output /*mux_wire*/ logic[31:0] rdata,
	output /*mux_wire*/ logic[1:0] rresp,
	output /*mux_wire*/ logic rvalid,
	input wire rready,
	output /*state*/ logic[31:0] input_regs[3:0],
	output /*mux_wire*/ logic start,
	input wire finish,
	input wire[31:0] output_regs[5:0]
);

genvar _g0;
/*state*/ logic[31:0] stored_output_regs[5:0];
/*state*/ logic reg_ctrl_ap_idle;
/*state*/ logic reg_ctrl_ap_done;
/*mux_wire*/ logic reg_ctrl_ap_ready;
/*state*/ logic reg_ctrl_ap_start;
/*state*/ logic[9:0] stored_addr;
/*state*/ logic stored_addr_valid;
/*state*/ logic[1:0] last_bresp;
/*state*/ logic last_werr_valid;
wire _4;
assign _4 = !stored_addr_valid;
wire _6;
assign _6 = _4 & aresetn;
wire _9;
assign _9 = !last_werr_valid;
wire _10;
assign _10 = stored_addr_valid & _9;
wire _15;
assign _15 = awready & awvalid;
wire[9:0] _17;
assign _17 = awaddr / 3'd4;
wire _20;
assign _20 = wready & wvalid;
localparam[1:0] RESP_SLVERR = 2'b10;
wire _22;
assign _22 = stored_addr == 1'd0;
wire _23 = wstrb[0];
wire _24 = wdata[0];
wire _25;
assign _25 = _23 & _24;
localparam[1:0] RESP_OKAY = 2'b00;
wire _28;
assign _28 = stored_addr >= 3'd4;
wire _31;
assign _31 = stored_addr < 4'd8;
wire _32;
assign _32 = _28 & _31;
/*mux_wire*/ logic[1:0] write_idx;
/*mux_wire*/ logic[9:0] _IntNarrow_in;
wire[2:0] _IntNarrow_out;
wire[1:0] _34;
assign _34 = _IntNarrow_out - 3'd4;
wire _35 = wstrb[0];
wire[7:0] _37;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _37[_g0] = wdata[_g0];
end
endgenerate
wire _38 = wstrb[1];
wire[7:0] _40;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _40[_g0] = wdata[8 + _g0];
end
endgenerate
wire _41 = wstrb[2];
wire[7:0] _43;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _43[_g0] = wdata[16 + _g0];
end
endgenerate
wire _44 = wstrb[3];
wire[7:0] _46;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _46[_g0] = wdata[24 + _g0];
end
endgenerate
localparam[1:0] RESP_OKAY_2 = 2'b00;
wire _49;
assign _49 = bready & bvalid;
/*state*/ logic last_rdata_valid;
/*state*/ logic[31:0] last_rdata;
/*state*/ logic[1:0] last_rresp;
/*mux_wire*/ logic[31:0] regs_read_multiplexer[9:0];
wire _55;
assign _55 = !last_rdata_valid;
wire _57;
assign _57 = _55 & aresetn;
wire _61;
assign _61 = arready & arvalid;
localparam[1:0] RESP_SLVERR_2 = 2'b10;
/*mux_wire*/ logic[9:0] read_addr;
wire[9:0] _63;
assign _63 = araddr / 3'd4;
wire _65;
assign _65 = read_addr == 1'd0;
/*mux_wire*/ logic _Repeat_v;
wire[27:0] _Repeat_result;
localparam[1:0] RESP_OKAY_3 = 2'b00;
wire _72;
assign _72 = read_addr >= 3'd4;
wire _75;
assign _75 = read_addr < 4'd14;
wire _76;
assign _76 = _72 & _75;
/*mux_wire*/ logic[3:0] read_idx;
/*mux_wire*/ logic[9:0] _IntNarrow_2_in;
wire[3:0] _IntNarrow_2_out;
wire[3:0] _78;
assign _78 = _IntNarrow_2_out - 3'd4;
wire[31:0] _80 = regs_read_multiplexer[read_idx];
localparam[1:0] RESP_OKAY_4 = 2'b00;
wire _83;
assign _83 = rready & rvalid;
/*mux_wire*/ logic _cross_finish_in;
/*mux_wire*/ logic[31:0] _cross_finish_data_in[5:0];
wire _cross_finish_out;
wire[31:0] _cross_finish_data_out[5:0];
/*mux_wire*/ logic[31:0] output_regs_vs[5:0];
wire _89;
assign _89 = !aresetn;
/*mux_wire*/ logic _Repeat_2_v;
wire[31:0] _Repeat_2_result;
/*mux_wire*/ logic[31:0] _Repeat_3_v;
wire[31:0] _Repeat_3_result[3:0];
/*mux_wire*/ logic _Repeat_4_v;
wire[31:0] _Repeat_4_result;
/*mux_wire*/ logic[31:0] _Repeat_5_v;
wire[31:0] _Repeat_5_result[5:0];
IntNarrow_FROM_I_0_TO_I_1024_FROM_4_TO_8 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
Repeat_T_type_bool_SIZE_28 Repeat(
	.clk(aclk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
IntNarrow_FROM_I_0_TO_I_1024_FROM_4_TO_14 IntNarrow_2(
	.clk(aclk),
	.in(_IntNarrow_2_in),
	.out(_IntNarrow_2_out)
);
CrossAction_T_type_bool_32_6 cross_finish(
	.in_clk(aclk),
	.in(_cross_finish_in),
	.data_in(_cross_finish_data_in),
	.out(_cross_finish_out),
	.data_out(_cross_finish_data_out)
);
Repeat_T_type_bool_SIZE_32 Repeat_2(
	.clk(aclk),
	.v(_Repeat_2_v),
	.result(_Repeat_2_result)
);
Repeat_T_type_bool_32_SIZE_4 Repeat_3(
	.clk(aclk),
	.v(_Repeat_3_v),
	.result(_Repeat_3_result)
);
Repeat_T_type_bool_SIZE_32 Repeat_4(
	.clk(aclk),
	.v(_Repeat_4_v),
	.result(_Repeat_4_result)
);
Repeat_T_type_bool_32_SIZE_6 Repeat_5(
	.clk(aclk),
	.v(_Repeat_5_v),
	.result(_Repeat_5_result)
);
always_comb begin // combinatorial awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awready = 1'bx;
	awready = 1'b0;
	awready = _6;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awready = awready;
end
always_comb begin // combinatorial wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wready = 1'bx;
	wready = 1'b0;
	wready = _10;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wready = wready;
end
always_comb begin // combinatorial bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	bresp = 2'bxx;
	bresp = last_bresp;
end
always_comb begin // combinatorial bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	bvalid = 1'bx;
	bvalid = 1'b0;
	bvalid = last_werr_valid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	bvalid = bvalid;
end
always_comb begin // combinatorial arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arready = 1'bx;
	arready = 1'b0;
	arready = _57;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arready = arready;
end
always_comb begin // combinatorial rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	rdata = last_rdata;
end
always_comb begin // combinatorial rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rresp = 2'bxx;
	rresp = last_rresp;
end
always_comb begin // combinatorial rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rvalid = 1'bx;
	rvalid = 1'b0;
	rvalid = last_rdata_valid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rvalid = rvalid;
end
always_ff @(posedge aclk) begin // state stored_output_regs
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
if(_cross_finish_out) stored_output_regs[_v0] <= output_regs_vs[_v0];
end
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
if(_89) stored_output_regs[_v0] <= _Repeat_5_result[_v0];
end
end
always_ff @(posedge aclk) begin // state input_regs
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_20) if(_32) if(_35) input_regs[write_idx][_v0] <= _37[_v0];
end
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_20) if(_32) if(_38) input_regs[write_idx][8 + _v0] <= _40[_v0];
end
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_20) if(_32) if(_41) input_regs[write_idx][16 + _v0] <= _43[_v0];
end
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_20) if(_32) if(_44) input_regs[write_idx][24 + _v0] <= _46[_v0];
end
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
if(_89) input_regs[_v0] <= _Repeat_3_result[_v0];
end
end
always_comb begin // combinatorial start
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	start = 1'bx;
	start = 1'b0;
	if(_20) if(_22) if(_25) start = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	start = start;
end
always_ff @(posedge aclk) begin // state reg_ctrl_ap_idle
	if(_20) if(_22) if(_25) reg_ctrl_ap_idle <= 1'b0;
	if(_61) if(_65) if(reg_ctrl_ap_done) reg_ctrl_ap_idle <= 1'b1;
	if(_cross_finish_out) reg_ctrl_ap_idle <= 1'b0;
	if(_89) reg_ctrl_ap_idle <= 1'b1;
end
always_ff @(posedge aclk) begin // state reg_ctrl_ap_done
	if(_61) if(_65) reg_ctrl_ap_done <= 1'b0;
	if(_cross_finish_out) reg_ctrl_ap_done <= 1'b1;
	if(_89) reg_ctrl_ap_done <= 1'b0;
end
always_comb begin // combinatorial reg_ctrl_ap_ready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	reg_ctrl_ap_ready = 1'bx;
	reg_ctrl_ap_ready = reg_ctrl_ap_done;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	reg_ctrl_ap_ready = reg_ctrl_ap_ready;
end
always_ff @(posedge aclk) begin // state reg_ctrl_ap_start
	if(_20) if(_22) if(_25) reg_ctrl_ap_start <= 1'b1;
	if(_cross_finish_out) reg_ctrl_ap_start <= 1'b0;
	if(_89) reg_ctrl_ap_start <= 1'b0;
end
always_ff @(posedge aclk) begin // state stored_addr
	if(_15) stored_addr <= _17;
end
always_ff @(posedge aclk) begin // state stored_addr_valid
	if(_15) stored_addr_valid <= 1'b1;
	if(_20) stored_addr_valid <= 1'b0;
	if(_89) stored_addr_valid <= 1'b0;
end
always_ff @(posedge aclk) begin // state last_bresp
	if(_20) last_bresp <= RESP_SLVERR;
	if(_20) if(_22) last_bresp <= RESP_OKAY;
	if(_20) if(_32) last_bresp <= RESP_OKAY_2;
end
always_ff @(posedge aclk) begin // state last_werr_valid
	if(_20) last_werr_valid <= 1'b1;
	if(_49) last_werr_valid <= 1'b0;
	if(_89) last_werr_valid <= 1'b0;
end
always_comb begin // combinatorial write_idx
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	write_idx = 2'dx;
	if(_20) if(_32) write_idx = _34;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 10'dx;
	if(_20) if(_32) _IntNarrow_in = stored_addr;
end
always_ff @(posedge aclk) begin // state last_rdata_valid
	if(_61) last_rdata_valid <= 1'b1;
	if(_83) last_rdata_valid <= 1'b0;
	if(_89) last_rdata_valid <= 1'b0;
end
always_ff @(posedge aclk) begin // state last_rdata
	if(_61) if(_65) last_rdata[0] <= reg_ctrl_ap_start;
	if(_61) if(_65) last_rdata[1] <= reg_ctrl_ap_done;
	if(_61) if(_65) last_rdata[2] <= reg_ctrl_ap_idle;
	if(_61) if(_65) last_rdata[3] <= reg_ctrl_ap_ready;
	for(int _v0 = 0; _v0 < 28; _v0 = _v0 + 1) begin
if(_61) if(_65) last_rdata[4 + _v0] <= _Repeat_result[_v0];
end
	if(_61) if(_76) last_rdata <= _80;
end
always_ff @(posedge aclk) begin // state last_rresp
	if(_61) last_rresp <= RESP_SLVERR_2;
	if(_61) if(_65) last_rresp <= RESP_OKAY_3;
	if(_61) if(_76) last_rresp <= RESP_OKAY_4;
end
always_comb begin // combinatorial regs_read_multiplexer
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	regs_read_multiplexer = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
regs_read_multiplexer[_v0] = input_regs[_v0];
end
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
regs_read_multiplexer[4 + _v0] = stored_output_regs[_v0];
end
end
always_comb begin // combinatorial read_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	read_addr = 10'dx;
	if(_61) read_addr = _63;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	if(_61) if(_65) _Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
always_comb begin // combinatorial read_idx
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	read_idx = 4'dx;
	if(_61) if(_76) read_idx = _78;
end
always_comb begin // combinatorial _IntNarrow_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_2_in = 10'dx;
	if(_61) if(_76) _IntNarrow_2_in = read_addr;
end
always_comb begin // combinatorial _cross_finish_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_finish_in = 1'bx;
	_cross_finish_in = 1'b0;
	if(finish) _cross_finish_in = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_finish_in = _cross_finish_in;
end
always_comb begin // combinatorial _cross_finish_data_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_finish_data_in = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
if(finish) _cross_finish_data_in[_v0] = output_regs[_v0];
end
end
always_comb begin // combinatorial output_regs_vs
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	output_regs_vs = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
if(_cross_finish_out) output_regs_vs[_v0] = _cross_finish_data_out[_v0];
end
end
always_comb begin // combinatorial _Repeat_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_2_v = 1'bx;
	if(_89) _Repeat_2_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_2_v = _Repeat_2_v;
end
always_comb begin // combinatorial _Repeat_3_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_3_v = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_89) _Repeat_3_v = _Repeat_2_result;
end
always_comb begin // combinatorial _Repeat_4_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_4_v = 1'bx;
	if(_89) _Repeat_4_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_4_v = _Repeat_4_v;
end
always_comb begin // combinatorial _Repeat_5_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_5_v = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_89) _Repeat_5_v = _Repeat_4_result;
end
endmodule

// Repeat #(T: type bool #()[32], SIZE: 6)
module Repeat_T_type_bool_32_SIZE_6(
	input clk,
	input wire[31:0] v,
	output /*mux_wire*/ logic[31:0] result[5:0]
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
	result[4] = v;
	result[5] = v;
end
endmodule

// Repeat #(T: type bool #()[32], SIZE: 4)
module Repeat_T_type_bool_32_SIZE_4(
	input clk,
	input wire[31:0] v,
	output /*mux_wire*/ logic[31:0] result[3:0]
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
end
endmodule

// CrossAction #(T: type bool #()[32][6])
module CrossAction_T_type_bool_32_6(
	input in_clk,
	input wire in,
	input wire[31:0] data_in[5:0],
	output /*mux_wire*/ logic out,
	output /*mux_wire*/ logic[31:0] data_out[5:0]
);

/*mux_wire*/ logic _cross_valid_in;
/*mux_wire*/ logic[31:0] _cross_data_in[5:0];
wire _cross_valid_out;
wire[31:0] _cross_data_out[5:0];
CrossDomain_T_type_bool cross_valid(
	.in_clk(in_clk),
	.in(_cross_valid_in),
	.out(_cross_valid_out)
);
CrossDomain_T_type_bool_32_6 cross_data(
	.in_clk(in_clk),
	.in(_cross_data_in),
	.out(_cross_data_out)
);
always_comb begin // combinatorial _cross_valid_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_valid_in = 1'bx;
	if(in) _cross_valid_in = 1'b1;
	if(!in) _cross_valid_in = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_valid_in = _cross_valid_in;
end
always_comb begin // combinatorial _cross_data_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_data_in = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
if(in) _cross_data_in[_v0] = data_in[_v0];
end
end
always_comb begin // combinatorial out
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	out = 1'bx;
	out = 1'b0;
	if(_cross_valid_out) out = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	out = out;
end
always_comb begin // combinatorial data_out
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	data_out = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
if(_cross_valid_out) data_out[_v0] = _cross_data_out[_v0];
end
end
endmodule

// CrossDomain #(T: type bool #()[32][6])
module CrossDomain_T_type_bool_32_6(
	input in_clk,
	input wire[31:0] in[5:0],
	output /*mux_wire*/ logic[31:0] out[5:0]
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 1024, FROM: 4, TO: 14)
module IntNarrow_FROM_I_0_TO_I_1024_FROM_4_TO_14(
	input clk,
	input wire[9:0] in,
	output /*mux_wire*/ logic[3:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 1024, FROM: 4, TO: 8)
module IntNarrow_FROM_I_0_TO_I_1024_FROM_4_TO_8(
	input clk,
	input wire[9:0] in,
	output /*mux_wire*/ logic[2:0] out
);

	assign out = in;
endmodule

// test_burst_reader #()
module test_burst_reader(
	input clk
);

axi_array_burst_reader_AXI_WIDTH_64_ADDR_ALIGN_2_COUNT_TO_65536_ATO_18446744073709551616 reader(
	.aclk(clk),
	.aresetn(),
	.arvalid(),
	.arready(),
	.araddr(),
	.arlen(),
	.arsize(),
	.arburst(),
	.arprot(),
	.arcache(),
	.arqos(),
	.arlock(),
	.arregion(),
	.rvalid(),
	.rready(),
	.rdata(),
	.rresp(),
	.rlast(),
	.is_ready_to_receive_lots_of_data(),
	.element_packet_valid(),
	.elements(),
	.chunk_offset(),
	.chunk_length(),
	.last(),
	.max_in_flight(),
	.may_request_new_burst(),
	.request_new_burst(),
	.start_addr(),
	.count()
);
axi_realigning_burst_reader_T_type_bool_32_17_AXI_WIDTH_512_ADDR_ALIGN_4_COUNT_TO_65536_ATO_18446744073709551616 unalignedBigSingleObjectReader(
	.aclk(clk),
	.aresetn(),
	.arvalid(),
	.arready(),
	.araddr(),
	.arlen(),
	.arsize(),
	.arburst(),
	.arprot(),
	.arcache(),
	.arqos(),
	.arlock(),
	.arregion(),
	.rvalid(),
	.rready(),
	.rdata(),
	.rresp(),
	.rlast(),
	.max_in_flight(),
	.may_request_new_burst(),
	.request_new_burst(),
	.start_addr(),
	.count(),
	.is_ready_to_receive_lots_of_data(),
	.value_valid(),
	.value(),
	.last()
);
axi_realigning_burst_reader_T_type_bool_32_16_AXI_WIDTH_512_ADDR_ALIGN_64_COUNT_TO_65536_ATO_18446744073709551616 alignedBigSingleObjectReader(
	.aclk(clk),
	.aresetn(),
	.arvalid(),
	.arready(),
	.araddr(),
	.arlen(),
	.arsize(),
	.arburst(),
	.arprot(),
	.arcache(),
	.arqos(),
	.arlock(),
	.arregion(),
	.rvalid(),
	.rready(),
	.rdata(),
	.rresp(),
	.rlast(),
	.max_in_flight(),
	.may_request_new_burst(),
	.request_new_burst(),
	.start_addr(),
	.count(),
	.is_ready_to_receive_lots_of_data(),
	.value_valid(),
	.value(),
	.last()
);
endmodule

// axi_realigning_burst_reader #(T: type bool #()[32][16], AXI_WIDTH: 512, ADDR_ALIGN: 64, COUNT_TO: 65536, ATO: 18446744073709551616)
module axi_realigning_burst_reader_T_type_bool_32_16_AXI_WIDTH_512_ADDR_ALIGN_64_COUNT_TO_65536_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic arvalid,
	input wire arready,
	output /*mux_wire*/ logic[63:0] araddr,
	output /*mux_wire*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[511:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[15:0] count,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic value_valid,
	output /*mux_wire*/ logic[31:0] value[15:0],
	output /*mux_wire*/ logic last
);

/*mux_wire*/ logic _parent_aresetn;
wire _parent_arvalid;
wire[63:0] _parent_araddr;
wire[7:0] _parent_arlen;
wire[2:0] _parent_arsize;
wire[1:0] _parent_arburst;
wire[2:0] _parent_arprot;
wire[3:0] _parent_arcache;
wire[3:0] _parent_arqos;
wire _parent_arlock;
wire[3:0] _parent_arregion;
wire _parent_rready;
/*mux_wire*/ logic _parent_arready;
/*mux_wire*/ logic _parent_rvalid;
/*mux_wire*/ logic[511:0] _parent_rdata;
/*mux_wire*/ logic[1:0] _parent_rresp;
/*mux_wire*/ logic _parent_rlast;
/*mux_wire*/ logic[10:0] _parent_max_in_flight;
wire _parent_may_request_new_burst;
wire[15:0] _22;
assign _22 = count * 1'd1;
/*mux_wire*/ logic _parent_request_new_burst;
/*mux_wire*/ logic[63:0] _parent_start_addr;
/*mux_wire*/ logic[15:0] _parent_count;
/*mux_wire*/ logic _parent_is_ready_to_receive_lots_of_data;
// (zero sized) stored_elements
// (zero sized) cur_element_store_align
wire _parent_element_packet_valid;
wire[511:0] _parent_elements[0:0];
// (zero sized) _parent_chunk_offset
wire[0:0] _parent_chunk_length;
wire _parent_last;
/*mux_wire*/ logic[511:0] elements[0:0];
// (zero sized) chunk_offset
/*mux_wire*/ logic[0:0] chunk_length;
/*mux_wire*/ logic last_2;
/*mux_wire*/ logic[511:0] elements_extended[0:0];
/*mux_wire*/ logic[511:0] rotated_elements[0:0];
// (zero sized) _31
// (zero sized) _32
/*mux_wire*/ logic[511:0] _RotateRight_data[0:0];
// (zero sized) _RotateRight_offset
wire[511:0] _RotateRight_rotated_data[0:0];
/*mux_wire*/ logic[0:0] rotated_strobe;
// (zero sized) _MakeStrobe_chunk_offset
/*mux_wire*/ logic[0:0] _MakeStrobe_chunk_length;
wire[0:0] _MakeStrobe_strobe;
/*mux_wire*/ logic[0:0] end_of_element;
wire[0:0] _37;
assign _37 = 1'd0 + chunk_length;
wire _39;
assign _39 = end_of_element >= 1'd1;
/*mux_wire*/ logic[511:0] resulting_value_bits;
wire[511:0] _40 = rotated_elements[0];
/*mux_wire*/ logic[511:0] _FromBits_bits;
wire[31:0] _FromBits_value[15:0];
// (zero sized) _45
wire _47;
assign _47 = !aresetn;
axi_array_burst_reader_AXI_WIDTH_512_ADDR_ALIGN_64_COUNT_TO_65536_ATO_18446744073709551616 parent(
	.aclk(aclk),
	.aresetn(_parent_aresetn),
	.arvalid(_parent_arvalid),
	.arready(_parent_arready),
	.araddr(_parent_araddr),
	.arlen(_parent_arlen),
	.arsize(_parent_arsize),
	.arburst(_parent_arburst),
	.arprot(_parent_arprot),
	.arcache(_parent_arcache),
	.arqos(_parent_arqos),
	.arlock(_parent_arlock),
	.arregion(_parent_arregion),
	.rvalid(_parent_rvalid),
	.rready(_parent_rready),
	.rdata(_parent_rdata),
	.rresp(_parent_rresp),
	.rlast(_parent_rlast),
	.is_ready_to_receive_lots_of_data(_parent_is_ready_to_receive_lots_of_data),
	.element_packet_valid(_parent_element_packet_valid),
	.elements(_parent_elements),
	// (zero sized port) .chunk_offset(_parent_chunk_offset)
	.chunk_length(_parent_chunk_length),
	.last(_parent_last),
	.max_in_flight(_parent_max_in_flight),
	.may_request_new_burst(_parent_may_request_new_burst),
	.request_new_burst(_parent_request_new_burst),
	.start_addr(_parent_start_addr),
	.count(_parent_count)
);
RotateRight_T_type_bool_512_ARRAY_LEN_1 RotateRight(
	.clk(aclk),
	.data(_RotateRight_data),
	// (zero sized port) .offset(_RotateRight_offset)
	.rotated_data(_RotateRight_rotated_data)
);
MakeStrobe_STROBE_WIDTH_1 MakeStrobe(
	.clk(aclk),
	// (zero sized port) .chunk_offset(_MakeStrobe_chunk_offset)
	.chunk_length(_MakeStrobe_chunk_length),
	.strobe(_MakeStrobe_strobe)
);
FromBits_T_type_bool_32_16 FromBits(
	.clk(aclk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial _parent_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_aresetn = 1'bx;
	_parent_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_aresetn = _parent_aresetn;
end
always_comb begin // combinatorial arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arvalid = 1'bx;
	arvalid = _parent_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arvalid = arvalid;
end
always_comb begin // combinatorial araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	araddr = 64'dx;
	araddr = _parent_araddr;
end
always_comb begin // combinatorial arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlen = 8'dx;
	arlen = _parent_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = _parent_arsize;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _parent_arburst;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _parent_arprot;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _parent_arcache;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = _parent_arqos;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = _parent_arlock;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = _parent_arregion;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = _parent_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _parent_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_arready = 1'bx;
	_parent_arready = arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_arready = _parent_arready;
end
always_comb begin // combinatorial _parent_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rvalid = 1'bx;
	_parent_rvalid = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rvalid = _parent_rvalid;
end
always_comb begin // combinatorial _parent_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rdata = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_parent_rdata = rdata;
end
always_comb begin // combinatorial _parent_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rresp = 2'bxx;
	_parent_rresp = rresp;
end
always_comb begin // combinatorial _parent_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rlast = 1'bx;
	_parent_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rlast = _parent_rlast;
end
always_comb begin // combinatorial _parent_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_max_in_flight = 11'dx;
	_parent_max_in_flight = max_in_flight;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _parent_may_request_new_burst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial _parent_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_request_new_burst = 1'bx;
	_parent_request_new_burst = 1'b0;
	if(request_new_burst) _parent_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_request_new_burst = _parent_request_new_burst;
end
always_comb begin // combinatorial _parent_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_start_addr = 64'dx;
	if(request_new_burst) _parent_start_addr = start_addr;
end
always_comb begin // combinatorial _parent_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_count = 16'dx;
	if(request_new_burst) _parent_count = _22;
end
always_comb begin // combinatorial _parent_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_is_ready_to_receive_lots_of_data = 1'bx;
	_parent_is_ready_to_receive_lots_of_data = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_is_ready_to_receive_lots_of_data = _parent_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value_valid = 1'bx;
	value_valid = 1'b0;
	if(_parent_element_packet_valid) if(_39) value_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	value_valid = value_valid;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) value[_v0] = _FromBits_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_parent_element_packet_valid) if(_39) last = last_2;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements[_v0] = _parent_elements[_v0];
end
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 1'dx;
	if(_parent_element_packet_valid) chunk_length = _parent_chunk_length;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunk_length = chunk_length;
end
always_comb begin // combinatorial last_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last_2 = 1'bx;
	if(_parent_element_packet_valid) last_2 = _parent_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last_2 = last_2;
end
always_comb begin // combinatorial elements_extended
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_extended = '{512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements_extended[_v0] = elements[_v0];
end
end
always_comb begin // combinatorial rotated_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_elements = '{512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) rotated_elements[_v0] = _RotateRight_rotated_data[_v0];
end
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = '{512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) _RotateRight_data[_v0] = elements_extended[_v0];
end
end
always_comb begin // combinatorial rotated_strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_strobe = 1'bx;
	if(_parent_element_packet_valid) rotated_strobe = _MakeStrobe_strobe;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rotated_strobe = rotated_strobe;
end
always_comb begin // combinatorial _MakeStrobe_chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_length = 1'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_length = chunk_length;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_MakeStrobe_chunk_length = _MakeStrobe_chunk_length;
end
always_comb begin // combinatorial end_of_element
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	end_of_element = 1'dx;
	if(_parent_element_packet_valid) end_of_element = _37;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	end_of_element = end_of_element;
end
always_comb begin // combinatorial resulting_value_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	resulting_value_bits = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 512; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) resulting_value_bits[_v0] = _40[_v0];
end
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_parent_element_packet_valid) if(_39) _FromBits_bits = resulting_value_bits;
end
endmodule

// FromBits #(T: type bool #()[32][16])
module FromBits_T_type_bool_32_16(
	input clk,
	input wire[511:0] bits,
	output /*mux_wire*/ logic[31:0] value[15:0]
);

genvar _g0;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign value[_g0] = bits[(_g0) * 32 +: 32];
end
endgenerate
endmodule

// MakeStrobe #(STROBE_WIDTH: 1)
module MakeStrobe_STROBE_WIDTH_1(
	input clk,
	// (zero sized) input chunk_offset
	input wire[0:0] chunk_length,
	output /*mux_wire*/ logic[0:0] strobe
);

/*mux_wire*/ logic[0:0] chunk_bits;
wire _2;
assign _2 = chunk_length > 1'd0;
/*mux_wire*/ logic[0:0] _RotateRight_data;
// (zero sized) _RotateRight_offset
wire[0:0] _RotateRight_rotated_data;
RotateRight_T_type_bool_ARRAY_LEN_1 RotateRight(
	.clk(clk),
	.data(_RotateRight_data),
	// (zero sized port) .offset(_RotateRight_offset)
	.rotated_data(_RotateRight_rotated_data)
);
always_comb begin // combinatorial strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	strobe = 1'bx;
	strobe = _RotateRight_rotated_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	strobe = strobe;
end
always_comb begin // combinatorial chunk_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_bits = 1'bx;
	if(_2) chunk_bits[0] = 1'b1;
	if(!_2) chunk_bits[0] = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunk_bits = chunk_bits;
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = 1'bx;
	_RotateRight_data = chunk_bits;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_RotateRight_data = _RotateRight_data;
end
endmodule

// RotateRight #(T: type bool #(), ARRAY_LEN: 1)
module RotateRight_T_type_bool_ARRAY_LEN_1(
	input clk,
	input wire[0:0] data,
	// (zero sized) input offset
	output /*mux_wire*/ logic[0:0] rotated_data
);

// (zero sized) offset_bits
// (zero sized) _UIntToBits_value
// (zero sized) _UIntToBits_bits
/*mux_wire*/ logic[0:0] rotate_stages[0:0];
wire[0:0] _3 = rotate_stages[0];
UIntToBits_NUM_BITS_0 UIntToBits(
	.clk(clk)
	// (zero sized port) .value(_UIntToBits_value)
	// (zero sized port) .bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = 1'bx;
	rotated_data = _3;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rotated_data = rotated_data;
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{1'bx};
	rotate_stages[0] = data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rotate_stages = rotate_stages;
end
endmodule

// RotateRight #(T: type bool #()[512], ARRAY_LEN: 1)
module RotateRight_T_type_bool_512_ARRAY_LEN_1(
	input clk,
	input wire[511:0] data[0:0],
	// (zero sized) input offset
	output /*mux_wire*/ logic[511:0] rotated_data[0:0]
);

genvar _g0;
// (zero sized) offset_bits
// (zero sized) _UIntToBits_value
// (zero sized) _UIntToBits_bits
/*mux_wire*/ logic[511:0] rotate_stages[0:0][0:0];
wire[511:0] _3[0:0];
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _3[_g0] = rotate_stages[0][_g0];
end
endgenerate
UIntToBits_NUM_BITS_0 UIntToBits(
	.clk(clk)
	// (zero sized port) .value(_UIntToBits_value)
	// (zero sized port) .bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = '{512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
rotated_data[_v0] = _3[_v0];
end
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{'{512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
rotate_stages[0][_v0] = data[_v0];
end
end
endmodule

// axi_array_burst_reader #(AXI_WIDTH: 512, ADDR_ALIGN: 64, COUNT_TO: 65536, ATO: 18446744073709551616)
module axi_array_burst_reader_AXI_WIDTH_512_ADDR_ALIGN_64_COUNT_TO_65536_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*state*/ logic arvalid,
	input wire arready,
	output /*state*/ logic[63:0] araddr,
	output /*state*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[511:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic element_packet_valid,
	output /*mux_wire*/ logic[511:0] elements[0:0],
	// (zero sized) output chunk_offset
	output /*mux_wire*/ logic[0:0] chunk_length,
	output /*mux_wire*/ logic last,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[15:0] count
);

/*latency*/ logic _arvalid_D1; always_ff @(posedge aclk) begin _arvalid_D1 <= arvalid; end
/*latency*/ logic _request_new_burst_D1; always_ff @(posedge aclk) begin _request_new_burst_D1 <= request_new_burst; end
genvar _g0;
localparam[1:0] _1 = 2'b01;
localparam[2:0] _2 = 3'b000;
localparam[3:0] _3 = 4'b0010;
/*mux_wire*/ logic[1:0] _rresp;
/*mux_wire*/ logic _rlast;
/*state*/ logic[11:0] num_in_flight;
/*state*/ logic last_burst_in_flight;
/*mux_wire*/ logic[63:0] next_araddr;
/*latency*/ logic[63:0] _next_araddr_D0; always_ff @(posedge aclk) begin _next_araddr_D0 <= next_araddr; end
wire[57:0] _cur_start_chunk_addr_old;
/*mux_wire*/ logic[57:0] _BitwiseIntConcat_upper;
/*mux_wire*/ logic[5:0] _BitwiseIntConcat_lower;
wire[63:0] _BitwiseIntConcat_v;
/*mux_wire*/ logic[5:0] next_arlen;
/*mux_wire*/ logic next_last_burst_in_flight;
/*latency*/ logic _next_last_burst_in_flight_D0; always_ff @(posedge aclk) begin _next_last_burst_in_flight_D0 <= next_last_burst_in_flight; end
/*mux_wire*/ logic[51:0] cur_burst_addr;
/*mux_wire*/ logic[5:0] cur_align;
/*mux_wire*/ logic[57:0] _BitwiseIntSplit_v;
wire[51:0] _BitwiseIntSplit_upper;
wire[5:0] _BitwiseIntSplit_lower;
/*mux_wire*/ logic chunks_are_left;
/*latency*/ logic _chunks_are_left_D0; always_ff @(posedge aclk) begin _chunks_are_left_D0 <= chunks_are_left; end
wire[16:0] _num_chunks_left_old;
/*latency*/ logic[16:0] __num_chunks_left_old_N1; always_ff @(posedge aclk) begin __num_chunks_left_old_N1 <= _num_chunks_left_old; end
/*latency*/ logic[16:0] __num_chunks_left_old_D0; always_ff @(posedge aclk) begin __num_chunks_left_old_D0 <= __num_chunks_left_old_N1; end
wire _14;
assign _14 = _num_chunks_left_old > 1'd0;
/*latency*/ logic __14_N1; always_ff @(posedge aclk) begin __14_N1 <= _14; end
/*mux_wire*/ logic[5:0] max_chunks_in_this_burst;
/*latency*/ logic[5:0] _max_chunks_in_this_burst_D0; always_ff @(posedge aclk) begin _max_chunks_in_this_burst_D0 <= max_chunks_in_this_burst; end
wire[5:0] _18;
assign _18 = 6'd63 - cur_align;
wire[6:0] _22;
assign _22 = max_chunks_in_this_burst + 1'd1;
wire _23;
assign _23 = __num_chunks_left_old_N1 <= _22;
/*latency*/ logic __23_D0; always_ff @(posedge aclk) begin __23_D0 <= _23; end
/*mux_wire*/ logic[16:0] _IntNarrow_in;
wire[6:0] _IntNarrow_out;
wire[5:0] _26;
assign _26 = _IntNarrow_out - 1'd1;
/*latency*/ logic[5:0] __26_D0; always_ff @(posedge aclk) begin __26_D0 <= _26; end
/*mux_wire*/ logic may_next_arvalid;
/*latency*/ logic _may_next_arvalid_D1; always_ff @(posedge aclk) begin _may_next_arvalid_D1 <= may_next_arvalid; end
wire _num_chunks_left_may_update;
wire _30;
assign _30 = _chunks_are_left_D0 & _num_chunks_left_may_update;
wire _cur_start_chunk_addr_may_update;
wire _32;
assign _32 = _30 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
wire _34;
assign _34 = _32 & _LatencyOffset_out;
wire signed[11:0] _37;
assign _37 = max_in_flight - 7'd64;
wire _38;
assign _38 = $signed({1'b0, num_in_flight}) <= _37;
wire _39;
assign _39 = _34 & _38;
/*mux_wire*/ logic[52:0] next_burst_addr;
wire[52:0] _45;
assign _45 = cur_burst_addr + 1'd1;
/*latency*/ logic[52:0] __45_D0; always_ff @(posedge aclk) begin __45_D0 <= _45; end
/*latency*/ logic[52:0] __45_D1; always_ff @(posedge aclk) begin __45_D1 <= __45_D0; end
/*mux_wire*/ logic[52:0] _BitwiseIntConcat_2_upper;
/*mux_wire*/ logic[5:0] _BitwiseIntConcat_2_lower;
wire[58:0] _BitwiseIntConcat_2_v;
/*mux_wire*/ logic[58:0] _IntNarrow_2_in;
wire[57:0] _IntNarrow_2_out;
/*mux_wire*/ logic _cur_start_chunk_addr_update;
/*mux_wire*/ logic[57:0] _cur_start_chunk_addr_new;
/*mux_wire*/ logic[16:0] next_num_chunks_left;
wire[6:0] _53;
assign _53 = next_arlen + 1'd1;
wire signed[17:0] _54;
assign _54 = __num_chunks_left_old_D0 - _53;
/*mux_wire*/ logic signed[17:0] _IntNarrow_3_in;
wire[16:0] _IntNarrow_3_out;
/*mux_wire*/ logic _num_chunks_left_update;
/*mux_wire*/ logic[16:0] _num_chunks_left_new;
/*mux_wire*/ logic _BoolToInt_i;
wire[0:0] _BoolToInt_o;
wire signed[12:0] _64;
assign _64 = num_in_flight - _BoolToInt_o;
wire _66;
assign _66 = !arvalid;
wire _68;
assign _68 = _66 & may_next_arvalid;
wire[6:0] _71;
assign _71 = next_arlen + 1'd1;
/*mux_wire*/ logic _Ternary_cond;
/*mux_wire*/ logic[6:0] _Ternary_a;
/*mux_wire*/ logic[6:0] _Ternary_b;
wire[6:0] _Ternary_o;
wire signed[12:0] _73;
assign _73 = _64 + $signed({1'b0, _Ternary_o});
/*mux_wire*/ logic signed[12:0] _IntNarrow_4_in;
wire[11:0] _IntNarrow_4_out;
/*state*/ logic[0:0] final_chunk_align;
// (zero sized) cur_chunk_align
/*mux_wire*/ logic[511:0] elements_2[0:0];
wire[511:0] _75;
generate
for(_g0 = 0; _g0 < 512; _g0 = _g0 + 1) begin
assign _75[_g0] = rdata[_g0];
end
endgenerate
/*mux_wire*/ logic[0:0] num_chunk_elements;
/*mux_wire*/ logic is_last;
wire _78;
assign _78 = num_in_flight == 1'd1;
wire _80;
assign _80 = _78 & last_burst_in_flight;
wire[0:0] _84;
assign _84 = final_chunk_align - 1'd0;
/*mux_wire*/ logic[0:0] _IntNarrow_5_in;
wire[0:0] _IntNarrow_5_out;
wire[0:0] _86;
assign _86 = 1'd1 - 1'd0;
wire _94;
assign _94 = !chunks_are_left;
/*latency*/ logic __94_D0; always_ff @(posedge aclk) begin __94_D0 <= _94; end
wire _96;
assign _96 = __94_D0 & _num_chunks_left_may_update;
wire _98;
assign _98 = _96 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic[57:0] chunk_addr;
/*latency*/ logic[57:0] _chunk_addr_D1; always_ff @(posedge aclk) begin _chunk_addr_D1 <= chunk_addr; end
// (zero sized) element_in_chunk_align
wire[57:0] _100;
assign _100 = start_addr / 7'd64;
/*mux_wire*/ logic[57:0] _BitwiseIntSplit_2_v;
wire[57:0] _BitwiseIntSplit_2_upper;
// (zero sized) _BitwiseIntSplit_2_lower
/*mux_wire*/ logic[15:0] chunk_count_bits;
// (zero sized) final_alignment
wire[15:0] _103;
assign _103 = count + 1'd0;
/*mux_wire*/ logic[15:0] _BitwiseIntSplit_3_v;
wire[15:0] _BitwiseIntSplit_3_upper;
// (zero sized) _BitwiseIntSplit_3_lower
/*mux_wire*/ logic[16:0] num_chunks;
/*mux_wire*/ logic is_no_chunks;
wire _106;
assign _106 = chunk_count_bits == 1'd0;
wire _112;
assign _112 = 1'd0 != 1'd0;
/*mux_wire*/ logic _BoolToInt_2_i;
wire[0:0] _BoolToInt_2_o;
wire[16:0] _113;
assign _113 = chunk_count_bits + _BoolToInt_2_o;
wire _119;
assign _119 = !is_no_chunks;
wire _122;
assign _122 = 1'd0 == 1'd0;
wire _123;
assign _123 = _119 & _122;
/*mux_wire*/ logic _BoolToInt_3_i;
wire[0:0] _BoolToInt_3_o;
/*mux_wire*/ logic[0:0] _BitwiseIntConcat_3_upper;
// (zero sized) _BitwiseIntConcat_3_lower
wire[0:0] _BitwiseIntConcat_3_v;
wire _127;
assign _127 = !aresetn;
/*mux_wire*/ logic _cur_start_chunk_addr_rst;
wire _129;
assign _129 = !aresetn;
/*mux_wire*/ logic _num_chunks_left_rst;
wire _131;
assign _131 = !aresetn;
SlowState_T_type_int_FROM_0_TO_288230376151711744_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1 cur_start_chunk_addr(
	.clk(aclk),
	.rst(_cur_start_chunk_addr_rst),
	.old(_cur_start_chunk_addr_old),
	.may_update(_cur_start_chunk_addr_may_update),
	.update(_cur_start_chunk_addr_update),
	.new_1(_cur_start_chunk_addr_new)
);
SlowState_T_type_int_FROM_0_TO_65539_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0 num_chunks_left(
	.clk(aclk),
	.rst(_num_chunks_left_rst),
	.old(_num_chunks_left_old),
	.may_update(_num_chunks_left_may_update),
	.update(_num_chunks_left_update),
	.new_1(_num_chunks_left_new)
);
BitwiseIntConcat_UPPER_TO_288230376151711744_LOWER_BITS_6 BitwiseIntConcat(
	.clk(aclk),
	.upper(_BitwiseIntConcat_upper),
	.lower(_BitwiseIntConcat_lower),
	.v(_BitwiseIntConcat_v)
);
BitwiseIntSplit_TO_288230376151711744_LOWER_BITS_6 BitwiseIntSplit(
	.clk(aclk),
	.v(_BitwiseIntSplit_v),
	.upper(_BitwiseIntSplit_upper),
	.lower(_BitwiseIntSplit_lower)
);
IntNarrow_FROM_I_0_TO_I_65539_FROM_1_TO_65 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
LatencyOffset_T_type_bool_OFFSET_192 LatencyOffset(
	.clk(aclk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
BitwiseIntConcat_UPPER_TO_4503599627370497_LOWER_BITS_6 BitwiseIntConcat_2(
	.clk(aclk),
	.upper(_BitwiseIntConcat_2_upper),
	.lower(_BitwiseIntConcat_2_lower),
	.v(_BitwiseIntConcat_2_v)
);
IntNarrow_FROM_I_0_TO_I_288230376151711808_FROM_0_TO_288230376151711744 IntNarrow_2(
	.clk(aclk),
	.in(_IntNarrow_2_in),
	.out(_IntNarrow_2_out)
);
IntNarrow_FROM_I_64_TO_I_65538_FROM_0_TO_65539 IntNarrow_3(
	.clk(aclk),
	.in(_IntNarrow_3_in),
	.out(_IntNarrow_3_out)
);
BoolToInt BoolToInt(
	.clk(aclk),
	.i(_BoolToInt_i),
	.o(_BoolToInt_o)
);
Ternary_T_type_int_FROM_0_TO_65 Ternary(
	.clk(aclk),
	.cond(_Ternary_cond),
	.a(_Ternary_a),
	.b(_Ternary_b),
	.o(_Ternary_o)
);
IntNarrow_FROM_I_1_TO_I_3256_FROM_0_TO_3192 IntNarrow_4(
	.clk(aclk),
	.in(_IntNarrow_4_in),
	.out(_IntNarrow_4_out)
);
IntNarrow_FROM_I_0_TO_I_2_FROM_0_TO_2 IntNarrow_5(
	.clk(aclk),
	.in(_IntNarrow_5_in),
	.out(_IntNarrow_5_out)
);
BitwiseIntSplit_TO_288230376151711744_LOWER_BITS_0 BitwiseIntSplit_2(
	.clk(aclk),
	.v(_BitwiseIntSplit_2_v),
	.upper(_BitwiseIntSplit_2_upper)
	// (zero sized port) .lower(_BitwiseIntSplit_2_lower)
);
BitwiseIntSplit_TO_65536_LOWER_BITS_0 BitwiseIntSplit_3(
	.clk(aclk),
	.v(_BitwiseIntSplit_3_v),
	.upper(_BitwiseIntSplit_3_upper)
	// (zero sized port) .lower(_BitwiseIntSplit_3_lower)
);
BoolToInt BoolToInt_2(
	.clk(aclk),
	.i(_BoolToInt_2_i),
	.o(_BoolToInt_2_o)
);
BoolToInt BoolToInt_3(
	.clk(aclk),
	.i(_BoolToInt_3_i),
	.o(_BoolToInt_3_o)
);
BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_0 BitwiseIntConcat_3(
	.clk(aclk),
	.upper(_BitwiseIntConcat_3_upper),
	// (zero sized port) .lower(_BitwiseIntConcat_3_lower)
	.v(_BitwiseIntConcat_3_v)
);
always_ff @(posedge aclk) begin // state arvalid
	if(arvalid) if(arready) arvalid <= 1'b0;
	if(!arvalid) if(may_next_arvalid) arvalid <= 1'b1;
	if(_131) arvalid <= 1'b0;
end
always_ff @(posedge aclk) begin // state araddr
	if(!arvalid) if(may_next_arvalid) araddr <= _next_araddr_D0;
end
always_ff @(posedge aclk) begin // state arlen
	if(!arvalid) if(may_next_arvalid) arlen <= next_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = 3'd6;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _1;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _2;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _3;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = 1'd0;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = 1'd0;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rresp = 2'bxx;
	_rresp = rresp;
end
always_comb begin // combinatorial _rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rlast = 1'bx;
	_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_rlast = _rlast;
end
always_comb begin // combinatorial element_packet_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_packet_valid = 1'bx;
	element_packet_valid = 1'b0;
	if(rvalid) element_packet_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	element_packet_valid = element_packet_valid;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(rvalid) elements[_v0] = elements_2[_v0];
end
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 1'dx;
	if(rvalid) chunk_length = num_chunk_elements;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunk_length = chunk_length;
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(rvalid) last = is_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state num_in_flight
	num_in_flight <= _IntNarrow_4_out;
	if(_131) num_in_flight <= 1'd0;
end
always_ff @(posedge aclk) begin // state last_burst_in_flight
	if(!arvalid) if(may_next_arvalid) last_burst_in_flight <= _next_last_burst_in_flight_D0;
end
always_comb begin // combinatorial next_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_araddr = 64'dx;
	next_araddr = _BitwiseIntConcat_v;
end
always_comb begin // combinatorial _BitwiseIntConcat_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_upper = 58'dx;
	_BitwiseIntConcat_upper = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial _BitwiseIntConcat_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_lower = 6'dx;
	_BitwiseIntConcat_lower = 1'd0;
end
always_comb begin // combinatorial next_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_arlen = 6'dx;
	if(_chunks_are_left_D0) if(__23_D0) next_arlen = __26_D0;
	if(_chunks_are_left_D0) if(!__23_D0) next_arlen = _max_chunks_in_this_burst_D0;
end
always_comb begin // combinatorial next_last_burst_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_last_burst_in_flight = 1'bx;
	next_last_burst_in_flight = 1'b0;
	if(chunks_are_left) if(_23) next_last_burst_in_flight = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	next_last_burst_in_flight = next_last_burst_in_flight;
end
always_comb begin // combinatorial cur_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_burst_addr = 52'dx;
	cur_burst_addr = _BitwiseIntSplit_upper;
end
always_comb begin // combinatorial cur_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_align = 6'dx;
	cur_align = _BitwiseIntSplit_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_v = 58'dx;
	_BitwiseIntSplit_v = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial chunks_are_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunks_are_left = 1'bx;
	chunks_are_left = __14_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunks_are_left = chunks_are_left;
end
always_comb begin // combinatorial max_chunks_in_this_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	max_chunks_in_this_burst = 6'dx;
	if(chunks_are_left) max_chunks_in_this_burst = _18;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 17'dx;
	if(chunks_are_left) if(_23) _IntNarrow_in = __num_chunks_left_old_N1;
end
always_comb begin // combinatorial may_next_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_next_arvalid = 1'bx;
	may_next_arvalid = _39;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_next_arvalid = may_next_arvalid;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial next_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_burst_addr = 53'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) next_burst_addr = __45_D1;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_upper = 53'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_upper = next_burst_addr;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_lower = 6'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_lower = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_2_in = 59'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _IntNarrow_2_in = _BitwiseIntConcat_2_v;
end
always_comb begin // combinatorial _cur_start_chunk_addr_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_update = 1'bx;
	_cur_start_chunk_addr_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _cur_start_chunk_addr_update = 1'b1;
	if(request_new_burst) _cur_start_chunk_addr_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_update = _cur_start_chunk_addr_update;
end
always_comb begin // combinatorial _cur_start_chunk_addr_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_new = 58'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _cur_start_chunk_addr_new = _IntNarrow_2_out;
	if(_request_new_burst_D1) _cur_start_chunk_addr_new = _chunk_addr_D1;
end
always_comb begin // combinatorial next_num_chunks_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_num_chunks_left = 17'dx;
	if(!arvalid) if(may_next_arvalid) next_num_chunks_left = _IntNarrow_3_out;
end
always_comb begin // combinatorial _IntNarrow_3_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_3_in = 18'sdx;
	if(!arvalid) if(may_next_arvalid) _IntNarrow_3_in = _54;
end
always_comb begin // combinatorial _num_chunks_left_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_update = 1'bx;
	_num_chunks_left_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_update = 1'b1;
	if(request_new_burst) _num_chunks_left_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_update = _num_chunks_left_update;
end
always_comb begin // combinatorial _num_chunks_left_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_new = 17'dx;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_new = next_num_chunks_left;
	if(request_new_burst) _num_chunks_left_new = num_chunks;
end
always_comb begin // combinatorial _BoolToInt_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_i = 1'bx;
	_BoolToInt_i = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_i = _BoolToInt_i;
end
always_comb begin // combinatorial _Ternary_cond
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_cond = 1'bx;
	_Ternary_cond = _68;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Ternary_cond = _Ternary_cond;
end
always_comb begin // combinatorial _Ternary_a
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_a = 7'dx;
	_Ternary_a = _71;
end
always_comb begin // combinatorial _Ternary_b
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_b = 7'dx;
	_Ternary_b = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_4_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_4_in = 13'sdx;
	_IntNarrow_4_in = _73;
end
always_ff @(posedge aclk) begin // state final_chunk_align
	if(request_new_burst) final_chunk_align <= _BitwiseIntConcat_3_v;
end
always_comb begin // combinatorial elements_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_2 = '{512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	if(rvalid) elements_2[0] = _75;
end
always_comb begin // combinatorial num_chunk_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunk_elements = 1'dx;
	if(rvalid) if(is_last) num_chunk_elements = _IntNarrow_5_out;
	if(rvalid) if(!is_last) num_chunk_elements = _86;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	num_chunk_elements = num_chunk_elements;
end
always_comb begin // combinatorial is_last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_last = 1'bx;
	if(rvalid) is_last = _80;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_last = is_last;
end
always_comb begin // combinatorial _IntNarrow_5_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_5_in = 1'dx;
	if(rvalid) if(is_last) _IntNarrow_5_in = _84;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_IntNarrow_5_in = _IntNarrow_5_in;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _98;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial chunk_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_addr = 58'dx;
	if(request_new_burst) chunk_addr = _BitwiseIntSplit_2_upper;
end
always_comb begin // combinatorial _BitwiseIntSplit_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_2_v = 58'dx;
	if(request_new_burst) _BitwiseIntSplit_2_v = _100;
end
always_comb begin // combinatorial chunk_count_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_count_bits = 16'dx;
	if(request_new_burst) chunk_count_bits = _BitwiseIntSplit_3_upper;
end
always_comb begin // combinatorial _BitwiseIntSplit_3_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_3_v = 16'dx;
	if(request_new_burst) _BitwiseIntSplit_3_v = _103;
end
always_comb begin // combinatorial num_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunks = 17'dx;
	if(request_new_burst) if(is_no_chunks) num_chunks = 1'd1;
	if(request_new_burst) if(!is_no_chunks) num_chunks = _113;
end
always_comb begin // combinatorial is_no_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_no_chunks = 1'bx;
	if(request_new_burst) is_no_chunks = _106;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_no_chunks = is_no_chunks;
end
always_comb begin // combinatorial _BoolToInt_2_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_2_i = 1'bx;
	if(request_new_burst) if(!is_no_chunks) _BoolToInt_2_i = _112;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_2_i = _BoolToInt_2_i;
end
always_comb begin // combinatorial _BoolToInt_3_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_3_i = 1'bx;
	if(request_new_burst) _BoolToInt_3_i = _123;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_3_i = _BoolToInt_3_i;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_upper = 1'dx;
	if(request_new_burst) _BitwiseIntConcat_3_upper = _BoolToInt_3_o;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BitwiseIntConcat_3_upper = _BitwiseIntConcat_3_upper;
end
always_comb begin // combinatorial _cur_start_chunk_addr_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_rst = 1'bx;
	_cur_start_chunk_addr_rst = _127;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_rst = _cur_start_chunk_addr_rst;
end
always_comb begin // combinatorial _num_chunks_left_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_rst = 1'bx;
	_num_chunks_left_rst = _129;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_rst = _num_chunks_left_rst;
end
endmodule

// BitwiseIntConcat #(UPPER_TO: 2, LOWER_BITS: 0)
module BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_0(
	input clk,
	input wire[0:0] upper,
	// (zero sized) input lower
	output /*mux_wire*/ logic[0:0] v
);

/*mux_wire*/ logic[0:0] v_bits;
// (zero sized) _UIntToBits_value
// (zero sized) _UIntToBits_bits
/*mux_wire*/ logic[0:0] _UIntToBits_2_value;
wire[0:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[0:0] _FromBits_bits;
wire[0:0] _FromBits_value;
UIntToBits_NUM_BITS_0 UIntToBits(
	.clk(clk)
	// (zero sized port) .value(_UIntToBits_value)
	// (zero sized port) .bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_1 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_2 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 1'dx;
	v = _FromBits_value;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	v = v;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 1'bx;
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_2_bits[_v0];
end
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	v_bits = v_bits;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 1'dx;
	_UIntToBits_2_value = upper;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_UIntToBits_2_value = _UIntToBits_2_value;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 1'bx;
	_FromBits_bits = v_bits;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_FromBits_bits = _FromBits_bits;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 2))
module FromBits_T_type_int_FROM_0_TO_2(
	input clk,
	input wire[0:0] bits,
	output /*mux_wire*/ logic[0:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 0)
module UIntToBits_NUM_BITS_0(
	input clk
	// (zero sized) input value
	// (zero sized) output bits
);

endmodule

// BitwiseIntSplit #(TO: 65536, LOWER_BITS: 0)
module BitwiseIntSplit_TO_65536_LOWER_BITS_0(
	input clk,
	input wire[15:0] v,
	output /*mux_wire*/ logic[15:0] upper
	// (zero sized) output lower
);

genvar _g0;
/*mux_wire*/ logic[15:0] v_bits;
/*mux_wire*/ logic[15:0] _UIntToBits_value;
wire[15:0] _UIntToBits_bits;
// (zero sized) _2
// (zero sized) _BitsToUInt_bits
// (zero sized) _BitsToUInt_value
wire[15:0] _3;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[15:0] _FromBits_bits;
wire[15:0] _FromBits_value;
UIntToBits_NUM_BITS_16 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_0 BitsToUInt(
	.clk(clk)
	// (zero sized port) .bits(_BitsToUInt_bits)
	// (zero sized port) .value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_65536 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 16'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 16'bxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 16'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 16'bxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 65536))
module FromBits_T_type_int_FROM_0_TO_65536(
	input clk,
	input wire[15:0] bits,
	output /*mux_wire*/ logic[15:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 16)
module UIntToBits_NUM_BITS_16(
	input clk,
	input wire[15:0] value,
	output /*mux_wire*/ logic[15:0] bits
);

	assign bits = value;
endmodule

// BitwiseIntSplit #(TO: 288230376151711744, LOWER_BITS: 0)
module BitwiseIntSplit_TO_288230376151711744_LOWER_BITS_0(
	input clk,
	input wire[57:0] v,
	output /*mux_wire*/ logic[57:0] upper
	// (zero sized) output lower
);

genvar _g0;
/*mux_wire*/ logic[57:0] v_bits;
/*mux_wire*/ logic[57:0] _UIntToBits_value;
wire[57:0] _UIntToBits_bits;
// (zero sized) _2
// (zero sized) _BitsToUInt_bits
// (zero sized) _BitsToUInt_value
wire[57:0] _3;
generate
for(_g0 = 0; _g0 < 58; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[57:0] _FromBits_bits;
wire[57:0] _FromBits_value;
UIntToBits_NUM_BITS_58 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_0 BitsToUInt(
	.clk(clk)
	// (zero sized port) .bits(_BitsToUInt_bits)
	// (zero sized port) .value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_288230376151711744 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 58'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 58'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 58'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 58'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// BitsToUInt #(NUM_BITS: 0)
module BitsToUInt_NUM_BITS_0(
	input clk
	// (zero sized) input bits
	// (zero sized) output value
);

endmodule

// IntNarrow #(FROM_I: 0, TO_I: 2, FROM: 0, TO: 2)
module IntNarrow_FROM_I_0_TO_I_2_FROM_0_TO_2(
	input clk,
	input wire[0:0] in,
	output /*mux_wire*/ logic[0:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: -64, TO_I: 65538, FROM: 0, TO: 65539)
module IntNarrow_FROM_I_64_TO_I_65538_FROM_0_TO_65539(
	input clk,
	input wire signed[17:0] in,
	output /*mux_wire*/ logic[16:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 65539, FROM: 1, TO: 65)
module IntNarrow_FROM_I_0_TO_I_65539_FROM_1_TO_65(
	input clk,
	input wire[16:0] in,
	output /*mux_wire*/ logic[6:0] out
);

	assign out = in;
endmodule

// SlowState #(T: type int #(FROM: 0, TO: 65539), RESET_TO: 0, OLD_DELAY: 2, NEW_DELAY: 0)
module SlowState_T_type_int_FROM_0_TO_65539_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0(
	input clk,
	input wire rst,
	output /*state*/ logic[16:0] old,
	output /*mux_wire*/ logic may_update,
	input wire update,
	input wire[16:0] new_1
);

genvar _g0;
/*mux_wire*/ logic _cross_rst_in;
/*mux_wire*/ logic[16:0] new_s;
/*mux_wire*/ logic update_s;
/*mux_wire*/ logic update_old;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
/*mux_wire*/ logic[16:0] new_old;
/*mux_wire*/ logic[16:0] _LatencyOffset_2_in;
wire[16:0] _LatencyOffset_2_out;
wire _cross_rst_out;
/*latency*/ logic __cross_rst_out_N1; always_ff @(posedge clk) begin __cross_rst_out_N1 <= _cross_rst_out; end
/*latency*/ logic __cross_rst_out_D0; always_ff @(posedge clk) begin __cross_rst_out_D0 <= __cross_rst_out_N1; end
/*state*/ logic[1:0] cooldown;
wire _8 = cooldown[0];
wire _11;
assign _11 = update_s | __cross_rst_out_D0;
/*mux_wire*/ logic _Repeat_v;
wire[1:0] _Repeat_result;
wire[0:0] _12;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _12[_g0] = cooldown[1 + _g0];
end
endgenerate
CrossDomain_T_type_bool cross_rst(
	.in_clk(clk),
	.in(_cross_rst_in),
	.out(_cross_rst_out)
);
LatencyOffset_T_type_bool_OFFSET_2 LatencyOffset(
	.clk(clk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
LatencyOffset_T_type_int_FROM_0_TO_65539_OFFSET_2 LatencyOffset_2(
	.clk(clk),
	.in(_LatencyOffset_2_in),
	.out(_LatencyOffset_2_out)
);
Repeat_T_type_bool_SIZE_2 Repeat(
	.clk(clk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
always_comb begin // combinatorial _cross_rst_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_rst_in = 1'bx;
	_cross_rst_in = rst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_rst_in = _cross_rst_in;
end
always_ff @(posedge clk) begin // state old
	if(_cross_rst_out) old <= 17'd0;
	if(!_cross_rst_out) if(update_old) old <= new_old;
end
always_comb begin // combinatorial new_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_s = 17'dx;
	if(update) new_s = new_1;
end
always_comb begin // combinatorial update_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_s = 1'bx;
	if(update) update_s = 1'b1;
	if(!update) update_s = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_s = update_s;
end
always_comb begin // combinatorial update_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_old = 1'bx;
	update_old = _LatencyOffset_out;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_old = update_old;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = update_s;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial new_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_old = 17'dx;
	new_old = _LatencyOffset_2_out;
end
always_comb begin // combinatorial _LatencyOffset_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_2_in = 17'dx;
	_LatencyOffset_2_in = new_s;
end
always_comb begin // combinatorial may_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_update = 1'bx;
	may_update = _8;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_update = may_update;
end
always_ff @(posedge clk) begin // state cooldown
	if(_11) cooldown <= _Repeat_result;
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(!_11) cooldown[_v0] <= _12[_v0];
end
	if(!_11) cooldown[1] <= 1'b1;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	if(_11) _Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
endmodule

// LatencyOffset #(T: type int #(FROM: 0, TO: 65539), OFFSET: -2)
module LatencyOffset_T_type_int_FROM_0_TO_65539_OFFSET_2(
	input clk,
	input wire[16:0] in,
	output /*mux_wire*/ logic[16:0] out
);

	assign out = in;
endmodule

// axi_realigning_burst_reader #(T: type bool #()[32][17], AXI_WIDTH: 512, ADDR_ALIGN: 4, COUNT_TO: 65536, ATO: 18446744073709551616)
module axi_realigning_burst_reader_T_type_bool_32_17_AXI_WIDTH_512_ADDR_ALIGN_4_COUNT_TO_65536_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic arvalid,
	input wire arready,
	output /*mux_wire*/ logic[63:0] araddr,
	output /*mux_wire*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[511:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[15:0] count,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic value_valid,
	output /*mux_wire*/ logic[31:0] value[16:0],
	output /*mux_wire*/ logic last
);

/*mux_wire*/ logic _parent_aresetn;
wire _parent_arvalid;
wire[63:0] _parent_araddr;
wire[7:0] _parent_arlen;
wire[2:0] _parent_arsize;
wire[1:0] _parent_arburst;
wire[2:0] _parent_arprot;
wire[3:0] _parent_arcache;
wire[3:0] _parent_arqos;
wire _parent_arlock;
wire[3:0] _parent_arregion;
wire _parent_rready;
/*mux_wire*/ logic _parent_arready;
/*mux_wire*/ logic _parent_rvalid;
/*mux_wire*/ logic[511:0] _parent_rdata;
/*mux_wire*/ logic[1:0] _parent_rresp;
/*mux_wire*/ logic _parent_rlast;
/*mux_wire*/ logic[10:0] _parent_max_in_flight;
wire _parent_may_request_new_burst;
wire[20:0] _22;
assign _22 = count * 5'd17;
/*mux_wire*/ logic _parent_request_new_burst;
/*mux_wire*/ logic[63:0] _parent_start_addr;
/*mux_wire*/ logic[20:0] _parent_count;
/*mux_wire*/ logic _parent_is_ready_to_receive_lots_of_data;
/*state*/ logic[31:0] stored_elements[15:0];
/*state*/ logic[4:0] cur_element_store_align;
wire _parent_element_packet_valid;
wire[31:0] _parent_elements[15:0];
wire[3:0] _parent_chunk_offset;
wire[4:0] _parent_chunk_length;
wire _parent_last;
/*mux_wire*/ logic[31:0] elements[15:0];
/*mux_wire*/ logic[3:0] chunk_offset;
/*mux_wire*/ logic[4:0] chunk_length;
/*mux_wire*/ logic last_2;
/*mux_wire*/ logic[31:0] elements_extended[16:0];
/*mux_wire*/ logic[31:0] rotated_elements[16:0];
wire signed[5:0] _31;
assign _31 = cur_element_store_align - chunk_offset;
wire[4:0] _32;
assign _32 = _31 + ((_31 < 0) ? 17 : 0); // == mod 17
/*mux_wire*/ logic[31:0] _RotateRight_data[16:0];
/*mux_wire*/ logic[4:0] _RotateRight_offset;
wire[31:0] _RotateRight_rotated_data[16:0];
/*mux_wire*/ logic[16:0] rotated_strobe;
/*mux_wire*/ logic[4:0] _MakeStrobe_chunk_offset;
/*mux_wire*/ logic[4:0] _MakeStrobe_chunk_length;
wire[16:0] _MakeStrobe_strobe;
/*mux_wire*/ logic[5:0] end_of_element;
wire[5:0] _37;
assign _37 = cur_element_store_align + chunk_length;
wire _39;
assign _39 = end_of_element >= 5'd17;
/*mux_wire*/ logic[543:0] resulting_value_bits;
wire[31:0] _40 = stored_elements[0];
wire _42;
assign _42 = cur_element_store_align > 1'd1;
wire[31:0] _43 = stored_elements[1];
wire[31:0] _44 = rotated_elements[1];
wire _46;
assign _46 = cur_element_store_align > 2'd2;
wire[31:0] _47 = stored_elements[2];
wire[31:0] _48 = rotated_elements[2];
wire _50;
assign _50 = cur_element_store_align > 2'd3;
wire[31:0] _51 = stored_elements[3];
wire[31:0] _52 = rotated_elements[3];
wire _54;
assign _54 = cur_element_store_align > 3'd4;
wire[31:0] _55 = stored_elements[4];
wire[31:0] _56 = rotated_elements[4];
wire _58;
assign _58 = cur_element_store_align > 3'd5;
wire[31:0] _59 = stored_elements[5];
wire[31:0] _60 = rotated_elements[5];
wire _62;
assign _62 = cur_element_store_align > 3'd6;
wire[31:0] _63 = stored_elements[6];
wire[31:0] _64 = rotated_elements[6];
wire _66;
assign _66 = cur_element_store_align > 3'd7;
wire[31:0] _67 = stored_elements[7];
wire[31:0] _68 = rotated_elements[7];
wire _70;
assign _70 = cur_element_store_align > 4'd8;
wire[31:0] _71 = stored_elements[8];
wire[31:0] _72 = rotated_elements[8];
wire _74;
assign _74 = cur_element_store_align > 4'd9;
wire[31:0] _75 = stored_elements[9];
wire[31:0] _76 = rotated_elements[9];
wire _78;
assign _78 = cur_element_store_align > 4'd10;
wire[31:0] _79 = stored_elements[10];
wire[31:0] _80 = rotated_elements[10];
wire _82;
assign _82 = cur_element_store_align > 4'd11;
wire[31:0] _83 = stored_elements[11];
wire[31:0] _84 = rotated_elements[11];
wire _86;
assign _86 = cur_element_store_align > 4'd12;
wire[31:0] _87 = stored_elements[12];
wire[31:0] _88 = rotated_elements[12];
wire _90;
assign _90 = cur_element_store_align > 4'd13;
wire[31:0] _91 = stored_elements[13];
wire[31:0] _92 = rotated_elements[13];
wire _94;
assign _94 = cur_element_store_align > 4'd14;
wire[31:0] _95 = stored_elements[14];
wire[31:0] _96 = rotated_elements[14];
wire _98;
assign _98 = cur_element_store_align > 4'd15;
wire[31:0] _99 = stored_elements[15];
wire[31:0] _100 = rotated_elements[15];
wire[31:0] _101 = rotated_elements[16];
/*mux_wire*/ logic[543:0] _FromBits_bits;
wire[31:0] _FromBits_value[16:0];
wire[4:0] _106;
assign _106 = end_of_element - ((end_of_element >= 17) ? 17 : 0); // == mod 17
wire _107 = rotated_strobe[0];
wire[31:0] _108 = rotated_elements[0];
wire _109 = rotated_strobe[1];
wire[31:0] _110 = rotated_elements[1];
wire _111 = rotated_strobe[2];
wire[31:0] _112 = rotated_elements[2];
wire _113 = rotated_strobe[3];
wire[31:0] _114 = rotated_elements[3];
wire _115 = rotated_strobe[4];
wire[31:0] _116 = rotated_elements[4];
wire _117 = rotated_strobe[5];
wire[31:0] _118 = rotated_elements[5];
wire _119 = rotated_strobe[6];
wire[31:0] _120 = rotated_elements[6];
wire _121 = rotated_strobe[7];
wire[31:0] _122 = rotated_elements[7];
wire _123 = rotated_strobe[8];
wire[31:0] _124 = rotated_elements[8];
wire _125 = rotated_strobe[9];
wire[31:0] _126 = rotated_elements[9];
wire _127 = rotated_strobe[10];
wire[31:0] _128 = rotated_elements[10];
wire _129 = rotated_strobe[11];
wire[31:0] _130 = rotated_elements[11];
wire _131 = rotated_strobe[12];
wire[31:0] _132 = rotated_elements[12];
wire _133 = rotated_strobe[13];
wire[31:0] _134 = rotated_elements[13];
wire _135 = rotated_strobe[14];
wire[31:0] _136 = rotated_elements[14];
wire _137 = rotated_strobe[15];
wire[31:0] _138 = rotated_elements[15];
wire _140;
assign _140 = !aresetn;
axi_array_burst_reader_AXI_WIDTH_512_ADDR_ALIGN_4_COUNT_TO_1114112_ATO_18446744073709551616 parent(
	.aclk(aclk),
	.aresetn(_parent_aresetn),
	.arvalid(_parent_arvalid),
	.arready(_parent_arready),
	.araddr(_parent_araddr),
	.arlen(_parent_arlen),
	.arsize(_parent_arsize),
	.arburst(_parent_arburst),
	.arprot(_parent_arprot),
	.arcache(_parent_arcache),
	.arqos(_parent_arqos),
	.arlock(_parent_arlock),
	.arregion(_parent_arregion),
	.rvalid(_parent_rvalid),
	.rready(_parent_rready),
	.rdata(_parent_rdata),
	.rresp(_parent_rresp),
	.rlast(_parent_rlast),
	.is_ready_to_receive_lots_of_data(_parent_is_ready_to_receive_lots_of_data),
	.element_packet_valid(_parent_element_packet_valid),
	.elements(_parent_elements),
	.chunk_offset(_parent_chunk_offset),
	.chunk_length(_parent_chunk_length),
	.last(_parent_last),
	.max_in_flight(_parent_max_in_flight),
	.may_request_new_burst(_parent_may_request_new_burst),
	.request_new_burst(_parent_request_new_burst),
	.start_addr(_parent_start_addr),
	.count(_parent_count)
);
RotateRight_T_type_bool_32_ARRAY_LEN_17 RotateRight(
	.clk(aclk),
	.data(_RotateRight_data),
	.offset(_RotateRight_offset),
	.rotated_data(_RotateRight_rotated_data)
);
MakeStrobe_STROBE_WIDTH_17 MakeStrobe(
	.clk(aclk),
	.chunk_offset(_MakeStrobe_chunk_offset),
	.chunk_length(_MakeStrobe_chunk_length),
	.strobe(_MakeStrobe_strobe)
);
FromBits_T_type_bool_32_17 FromBits(
	.clk(aclk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial _parent_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_aresetn = 1'bx;
	_parent_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_aresetn = _parent_aresetn;
end
always_comb begin // combinatorial arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arvalid = 1'bx;
	arvalid = _parent_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arvalid = arvalid;
end
always_comb begin // combinatorial araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	araddr = 64'dx;
	araddr = _parent_araddr;
end
always_comb begin // combinatorial arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlen = 8'dx;
	arlen = _parent_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = _parent_arsize;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _parent_arburst;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _parent_arprot;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _parent_arcache;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = _parent_arqos;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = _parent_arlock;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = _parent_arregion;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = _parent_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _parent_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_arready = 1'bx;
	_parent_arready = arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_arready = _parent_arready;
end
always_comb begin // combinatorial _parent_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rvalid = 1'bx;
	_parent_rvalid = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rvalid = _parent_rvalid;
end
always_comb begin // combinatorial _parent_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rdata = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_parent_rdata = rdata;
end
always_comb begin // combinatorial _parent_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rresp = 2'bxx;
	_parent_rresp = rresp;
end
always_comb begin // combinatorial _parent_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_rlast = 1'bx;
	_parent_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_rlast = _parent_rlast;
end
always_comb begin // combinatorial _parent_max_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_max_in_flight = 11'dx;
	_parent_max_in_flight = max_in_flight;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _parent_may_request_new_burst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial _parent_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_request_new_burst = 1'bx;
	_parent_request_new_burst = 1'b0;
	if(request_new_burst) _parent_request_new_burst = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_request_new_burst = _parent_request_new_burst;
end
always_comb begin // combinatorial _parent_start_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_start_addr = 64'dx;
	if(request_new_burst) _parent_start_addr = start_addr;
end
always_comb begin // combinatorial _parent_count
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_count = 21'dx;
	if(request_new_burst) _parent_count = _22;
end
always_comb begin // combinatorial _parent_is_ready_to_receive_lots_of_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_parent_is_ready_to_receive_lots_of_data = 1'bx;
	_parent_is_ready_to_receive_lots_of_data = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_parent_is_ready_to_receive_lots_of_data = _parent_is_ready_to_receive_lots_of_data;
end
always_comb begin // combinatorial value_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value_valid = 1'bx;
	value_valid = 1'b0;
	if(_parent_element_packet_valid) if(_39) value_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	value_valid = value_valid;
end
always_comb begin // combinatorial value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	value = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 17; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) value[_v0] = _FromBits_value[_v0];
end
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(_parent_element_packet_valid) if(_39) last = last_2;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state stored_elements
	if(_parent_element_packet_valid) if(_107) stored_elements[0] <= _108;
	if(_parent_element_packet_valid) if(_109) stored_elements[1] <= _110;
	if(_parent_element_packet_valid) if(_111) stored_elements[2] <= _112;
	if(_parent_element_packet_valid) if(_113) stored_elements[3] <= _114;
	if(_parent_element_packet_valid) if(_115) stored_elements[4] <= _116;
	if(_parent_element_packet_valid) if(_117) stored_elements[5] <= _118;
	if(_parent_element_packet_valid) if(_119) stored_elements[6] <= _120;
	if(_parent_element_packet_valid) if(_121) stored_elements[7] <= _122;
	if(_parent_element_packet_valid) if(_123) stored_elements[8] <= _124;
	if(_parent_element_packet_valid) if(_125) stored_elements[9] <= _126;
	if(_parent_element_packet_valid) if(_127) stored_elements[10] <= _128;
	if(_parent_element_packet_valid) if(_129) stored_elements[11] <= _130;
	if(_parent_element_packet_valid) if(_131) stored_elements[12] <= _132;
	if(_parent_element_packet_valid) if(_133) stored_elements[13] <= _134;
	if(_parent_element_packet_valid) if(_135) stored_elements[14] <= _136;
	if(_parent_element_packet_valid) if(_137) stored_elements[15] <= _138;
end
always_ff @(posedge aclk) begin // state cur_element_store_align
	if(_parent_element_packet_valid) cur_element_store_align <= _106;
	if(_140) cur_element_store_align <= 1'd0;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements[_v0] = _parent_elements[_v0];
end
end
always_comb begin // combinatorial chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_offset = 4'dx;
	if(_parent_element_packet_valid) chunk_offset = _parent_chunk_offset;
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 5'dx;
	if(_parent_element_packet_valid) chunk_length = _parent_chunk_length;
end
always_comb begin // combinatorial last_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last_2 = 1'bx;
	if(_parent_element_packet_valid) last_2 = _parent_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last_2 = last_2;
end
always_comb begin // combinatorial elements_extended
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_extended = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) elements_extended[_v0] = elements[_v0];
end
end
always_comb begin // combinatorial rotated_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 17; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) rotated_elements[_v0] = _RotateRight_rotated_data[_v0];
end
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 17; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) _RotateRight_data[_v0] = elements_extended[_v0];
end
end
always_comb begin // combinatorial _RotateRight_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_offset = 5'dx;
	if(_parent_element_packet_valid) _RotateRight_offset = _32;
end
always_comb begin // combinatorial rotated_strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_strobe = 17'bxxxxxxxxxxxxxxxxx;
	if(_parent_element_packet_valid) rotated_strobe = _MakeStrobe_strobe;
end
always_comb begin // combinatorial _MakeStrobe_chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_offset = 5'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_offset = cur_element_store_align;
end
always_comb begin // combinatorial _MakeStrobe_chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_MakeStrobe_chunk_length = 5'dx;
	if(_parent_element_packet_valid) _MakeStrobe_chunk_length = chunk_length;
end
always_comb begin // combinatorial end_of_element
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	end_of_element = 6'dx;
	if(_parent_element_packet_valid) end_of_element = _37;
end
always_comb begin // combinatorial resulting_value_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	resulting_value_bits = 544'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) resulting_value_bits[_v0] = _40[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_42) resulting_value_bits[32 + _v0] = _43[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_42) resulting_value_bits[32 + _v0] = _44[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_46) resulting_value_bits[64 + _v0] = _47[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_46) resulting_value_bits[64 + _v0] = _48[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_50) resulting_value_bits[96 + _v0] = _51[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_50) resulting_value_bits[96 + _v0] = _52[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_54) resulting_value_bits[128 + _v0] = _55[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_54) resulting_value_bits[128 + _v0] = _56[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_58) resulting_value_bits[160 + _v0] = _59[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_58) resulting_value_bits[160 + _v0] = _60[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_62) resulting_value_bits[192 + _v0] = _63[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_62) resulting_value_bits[192 + _v0] = _64[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_66) resulting_value_bits[224 + _v0] = _67[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_66) resulting_value_bits[224 + _v0] = _68[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_70) resulting_value_bits[256 + _v0] = _71[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_70) resulting_value_bits[256 + _v0] = _72[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_74) resulting_value_bits[288 + _v0] = _75[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_74) resulting_value_bits[288 + _v0] = _76[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_78) resulting_value_bits[320 + _v0] = _79[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_78) resulting_value_bits[320 + _v0] = _80[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_82) resulting_value_bits[352 + _v0] = _83[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_82) resulting_value_bits[352 + _v0] = _84[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_86) resulting_value_bits[384 + _v0] = _87[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_86) resulting_value_bits[384 + _v0] = _88[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_90) resulting_value_bits[416 + _v0] = _91[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_90) resulting_value_bits[416 + _v0] = _92[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_94) resulting_value_bits[448 + _v0] = _95[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_94) resulting_value_bits[448 + _v0] = _96[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(_98) resulting_value_bits[480 + _v0] = _99[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) if(!_98) resulting_value_bits[480 + _v0] = _100[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(_parent_element_packet_valid) if(_39) resulting_value_bits[512 + _v0] = _101[_v0];
end
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 544'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_parent_element_packet_valid) if(_39) _FromBits_bits = resulting_value_bits;
end
endmodule

// FromBits #(T: type bool #()[32][17])
module FromBits_T_type_bool_32_17(
	input clk,
	input wire[543:0] bits,
	output /*mux_wire*/ logic[31:0] value[16:0]
);

genvar _g0;
generate
for(_g0 = 0; _g0 < 17; _g0 = _g0 + 1) begin
assign value[_g0] = bits[(_g0) * 32 +: 32];
end
endgenerate
endmodule

// MakeStrobe #(STROBE_WIDTH: 17)
module MakeStrobe_STROBE_WIDTH_17(
	input clk,
	input wire[4:0] chunk_offset,
	input wire[4:0] chunk_length,
	output /*mux_wire*/ logic[16:0] strobe
);

/*mux_wire*/ logic[16:0] chunk_bits;
wire _2;
assign _2 = chunk_length > 1'd0;
wire _4;
assign _4 = chunk_length > 1'd1;
wire _6;
assign _6 = chunk_length > 2'd2;
wire _8;
assign _8 = chunk_length > 2'd3;
wire _10;
assign _10 = chunk_length > 3'd4;
wire _12;
assign _12 = chunk_length > 3'd5;
wire _14;
assign _14 = chunk_length > 3'd6;
wire _16;
assign _16 = chunk_length > 3'd7;
wire _18;
assign _18 = chunk_length > 4'd8;
wire _20;
assign _20 = chunk_length > 4'd9;
wire _22;
assign _22 = chunk_length > 4'd10;
wire _24;
assign _24 = chunk_length > 4'd11;
wire _26;
assign _26 = chunk_length > 4'd12;
wire _28;
assign _28 = chunk_length > 4'd13;
wire _30;
assign _30 = chunk_length > 4'd14;
wire _32;
assign _32 = chunk_length > 4'd15;
wire _34;
assign _34 = chunk_length > 5'd16;
/*mux_wire*/ logic[16:0] _RotateRight_data;
/*mux_wire*/ logic[4:0] _RotateRight_offset;
wire[16:0] _RotateRight_rotated_data;
RotateRight_T_type_bool_ARRAY_LEN_17 RotateRight(
	.clk(clk),
	.data(_RotateRight_data),
	.offset(_RotateRight_offset),
	.rotated_data(_RotateRight_rotated_data)
);
always_comb begin // combinatorial strobe
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	strobe = 17'bxxxxxxxxxxxxxxxxx;
	strobe = _RotateRight_rotated_data;
end
always_comb begin // combinatorial chunk_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_bits = 17'bxxxxxxxxxxxxxxxxx;
	if(_2) chunk_bits[0] = 1'b1;
	if(!_2) chunk_bits[0] = 1'b0;
	if(_4) chunk_bits[1] = 1'b1;
	if(!_4) chunk_bits[1] = 1'b0;
	if(_6) chunk_bits[2] = 1'b1;
	if(!_6) chunk_bits[2] = 1'b0;
	if(_8) chunk_bits[3] = 1'b1;
	if(!_8) chunk_bits[3] = 1'b0;
	if(_10) chunk_bits[4] = 1'b1;
	if(!_10) chunk_bits[4] = 1'b0;
	if(_12) chunk_bits[5] = 1'b1;
	if(!_12) chunk_bits[5] = 1'b0;
	if(_14) chunk_bits[6] = 1'b1;
	if(!_14) chunk_bits[6] = 1'b0;
	if(_16) chunk_bits[7] = 1'b1;
	if(!_16) chunk_bits[7] = 1'b0;
	if(_18) chunk_bits[8] = 1'b1;
	if(!_18) chunk_bits[8] = 1'b0;
	if(_20) chunk_bits[9] = 1'b1;
	if(!_20) chunk_bits[9] = 1'b0;
	if(_22) chunk_bits[10] = 1'b1;
	if(!_22) chunk_bits[10] = 1'b0;
	if(_24) chunk_bits[11] = 1'b1;
	if(!_24) chunk_bits[11] = 1'b0;
	if(_26) chunk_bits[12] = 1'b1;
	if(!_26) chunk_bits[12] = 1'b0;
	if(_28) chunk_bits[13] = 1'b1;
	if(!_28) chunk_bits[13] = 1'b0;
	if(_30) chunk_bits[14] = 1'b1;
	if(!_30) chunk_bits[14] = 1'b0;
	if(_32) chunk_bits[15] = 1'b1;
	if(!_32) chunk_bits[15] = 1'b0;
	if(_34) chunk_bits[16] = 1'b1;
	if(!_34) chunk_bits[16] = 1'b0;
end
always_comb begin // combinatorial _RotateRight_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_data = 17'bxxxxxxxxxxxxxxxxx;
	_RotateRight_data = chunk_bits;
end
always_comb begin // combinatorial _RotateRight_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_RotateRight_offset = 5'dx;
	_RotateRight_offset = chunk_offset;
end
endmodule

// RotateRight #(T: type bool #(), ARRAY_LEN: 17)
module RotateRight_T_type_bool_ARRAY_LEN_17(
	input clk,
	input wire[16:0] data,
	input wire[4:0] offset,
	output /*mux_wire*/ logic[16:0] rotated_data
);

/*mux_wire*/ logic[4:0] offset_bits;
/*mux_wire*/ logic[4:0] _UIntToBits_value;
wire[4:0] _UIntToBits_bits;
/*mux_wire*/ logic[16:0] rotate_stages[5:0];
/*mux_wire*/ logic[16:0] from;
wire[16:0] _3 = rotate_stages[0];
wire _4 = offset_bits[0];
wire _5 = from[16];
wire _6 = from[0];
wire _7 = offset_bits[0];
wire _8 = from[0];
wire _9 = from[1];
wire _10 = offset_bits[0];
wire _11 = from[1];
wire _12 = from[2];
wire _13 = offset_bits[0];
wire _14 = from[2];
wire _15 = from[3];
wire _16 = offset_bits[0];
wire _17 = from[3];
wire _18 = from[4];
wire _19 = offset_bits[0];
wire _20 = from[4];
wire _21 = from[5];
wire _22 = offset_bits[0];
wire _23 = from[5];
wire _24 = from[6];
wire _25 = offset_bits[0];
wire _26 = from[6];
wire _27 = from[7];
wire _28 = offset_bits[0];
wire _29 = from[7];
wire _30 = from[8];
wire _31 = offset_bits[0];
wire _32 = from[8];
wire _33 = from[9];
wire _34 = offset_bits[0];
wire _35 = from[9];
wire _36 = from[10];
wire _37 = offset_bits[0];
wire _38 = from[10];
wire _39 = from[11];
wire _40 = offset_bits[0];
wire _41 = from[11];
wire _42 = from[12];
wire _43 = offset_bits[0];
wire _44 = from[12];
wire _45 = from[13];
wire _46 = offset_bits[0];
wire _47 = from[13];
wire _48 = from[14];
wire _49 = offset_bits[0];
wire _50 = from[14];
wire _51 = from[15];
wire _52 = offset_bits[0];
wire _53 = from[15];
wire _54 = from[16];
/*mux_wire*/ logic[16:0] from_2;
wire[16:0] _55 = rotate_stages[1];
wire _56 = offset_bits[1];
wire _57 = from_2[15];
wire _58 = from_2[0];
wire _59 = offset_bits[1];
wire _60 = from_2[16];
wire _61 = from_2[1];
wire _62 = offset_bits[1];
wire _63 = from_2[0];
wire _64 = from_2[2];
wire _65 = offset_bits[1];
wire _66 = from_2[1];
wire _67 = from_2[3];
wire _68 = offset_bits[1];
wire _69 = from_2[2];
wire _70 = from_2[4];
wire _71 = offset_bits[1];
wire _72 = from_2[3];
wire _73 = from_2[5];
wire _74 = offset_bits[1];
wire _75 = from_2[4];
wire _76 = from_2[6];
wire _77 = offset_bits[1];
wire _78 = from_2[5];
wire _79 = from_2[7];
wire _80 = offset_bits[1];
wire _81 = from_2[6];
wire _82 = from_2[8];
wire _83 = offset_bits[1];
wire _84 = from_2[7];
wire _85 = from_2[9];
wire _86 = offset_bits[1];
wire _87 = from_2[8];
wire _88 = from_2[10];
wire _89 = offset_bits[1];
wire _90 = from_2[9];
wire _91 = from_2[11];
wire _92 = offset_bits[1];
wire _93 = from_2[10];
wire _94 = from_2[12];
wire _95 = offset_bits[1];
wire _96 = from_2[11];
wire _97 = from_2[13];
wire _98 = offset_bits[1];
wire _99 = from_2[12];
wire _100 = from_2[14];
wire _101 = offset_bits[1];
wire _102 = from_2[13];
wire _103 = from_2[15];
wire _104 = offset_bits[1];
wire _105 = from_2[14];
wire _106 = from_2[16];
/*mux_wire*/ logic[16:0] from_3;
wire[16:0] _107 = rotate_stages[2];
wire _108 = offset_bits[2];
wire _109 = from_3[13];
wire _110 = from_3[0];
wire _111 = offset_bits[2];
wire _112 = from_3[14];
wire _113 = from_3[1];
wire _114 = offset_bits[2];
wire _115 = from_3[15];
wire _116 = from_3[2];
wire _117 = offset_bits[2];
wire _118 = from_3[16];
wire _119 = from_3[3];
wire _120 = offset_bits[2];
wire _121 = from_3[0];
wire _122 = from_3[4];
wire _123 = offset_bits[2];
wire _124 = from_3[1];
wire _125 = from_3[5];
wire _126 = offset_bits[2];
wire _127 = from_3[2];
wire _128 = from_3[6];
wire _129 = offset_bits[2];
wire _130 = from_3[3];
wire _131 = from_3[7];
wire _132 = offset_bits[2];
wire _133 = from_3[4];
wire _134 = from_3[8];
wire _135 = offset_bits[2];
wire _136 = from_3[5];
wire _137 = from_3[9];
wire _138 = offset_bits[2];
wire _139 = from_3[6];
wire _140 = from_3[10];
wire _141 = offset_bits[2];
wire _142 = from_3[7];
wire _143 = from_3[11];
wire _144 = offset_bits[2];
wire _145 = from_3[8];
wire _146 = from_3[12];
wire _147 = offset_bits[2];
wire _148 = from_3[9];
wire _149 = from_3[13];
wire _150 = offset_bits[2];
wire _151 = from_3[10];
wire _152 = from_3[14];
wire _153 = offset_bits[2];
wire _154 = from_3[11];
wire _155 = from_3[15];
wire _156 = offset_bits[2];
wire _157 = from_3[12];
wire _158 = from_3[16];
/*mux_wire*/ logic[16:0] from_4;
wire[16:0] _159 = rotate_stages[3];
wire _160 = offset_bits[3];
wire _161 = from_4[9];
wire _162 = from_4[0];
wire _163 = offset_bits[3];
wire _164 = from_4[10];
wire _165 = from_4[1];
wire _166 = offset_bits[3];
wire _167 = from_4[11];
wire _168 = from_4[2];
wire _169 = offset_bits[3];
wire _170 = from_4[12];
wire _171 = from_4[3];
wire _172 = offset_bits[3];
wire _173 = from_4[13];
wire _174 = from_4[4];
wire _175 = offset_bits[3];
wire _176 = from_4[14];
wire _177 = from_4[5];
wire _178 = offset_bits[3];
wire _179 = from_4[15];
wire _180 = from_4[6];
wire _181 = offset_bits[3];
wire _182 = from_4[16];
wire _183 = from_4[7];
wire _184 = offset_bits[3];
wire _185 = from_4[0];
wire _186 = from_4[8];
wire _187 = offset_bits[3];
wire _188 = from_4[1];
wire _189 = from_4[9];
wire _190 = offset_bits[3];
wire _191 = from_4[2];
wire _192 = from_4[10];
wire _193 = offset_bits[3];
wire _194 = from_4[3];
wire _195 = from_4[11];
wire _196 = offset_bits[3];
wire _197 = from_4[4];
wire _198 = from_4[12];
wire _199 = offset_bits[3];
wire _200 = from_4[5];
wire _201 = from_4[13];
wire _202 = offset_bits[3];
wire _203 = from_4[6];
wire _204 = from_4[14];
wire _205 = offset_bits[3];
wire _206 = from_4[7];
wire _207 = from_4[15];
wire _208 = offset_bits[3];
wire _209 = from_4[8];
wire _210 = from_4[16];
/*mux_wire*/ logic[16:0] from_5;
wire[16:0] _211 = rotate_stages[4];
wire _212 = offset_bits[4];
wire _213 = from_5[1];
wire _214 = from_5[0];
wire _215 = offset_bits[4];
wire _216 = from_5[2];
wire _217 = from_5[1];
wire _218 = offset_bits[4];
wire _219 = from_5[3];
wire _220 = from_5[2];
wire _221 = offset_bits[4];
wire _222 = from_5[4];
wire _223 = from_5[3];
wire _224 = offset_bits[4];
wire _225 = from_5[5];
wire _226 = from_5[4];
wire _227 = offset_bits[4];
wire _228 = from_5[6];
wire _229 = from_5[5];
wire _230 = offset_bits[4];
wire _231 = from_5[7];
wire _232 = from_5[6];
wire _233 = offset_bits[4];
wire _234 = from_5[8];
wire _235 = from_5[7];
wire _236 = offset_bits[4];
wire _237 = from_5[9];
wire _238 = from_5[8];
wire _239 = offset_bits[4];
wire _240 = from_5[10];
wire _241 = from_5[9];
wire _242 = offset_bits[4];
wire _243 = from_5[11];
wire _244 = from_5[10];
wire _245 = offset_bits[4];
wire _246 = from_5[12];
wire _247 = from_5[11];
wire _248 = offset_bits[4];
wire _249 = from_5[13];
wire _250 = from_5[12];
wire _251 = offset_bits[4];
wire _252 = from_5[14];
wire _253 = from_5[13];
wire _254 = offset_bits[4];
wire _255 = from_5[15];
wire _256 = from_5[14];
wire _257 = offset_bits[4];
wire _258 = from_5[16];
wire _259 = from_5[15];
wire _260 = offset_bits[4];
wire _261 = from_5[0];
wire _262 = from_5[16];
wire[16:0] _263 = rotate_stages[5];
UIntToBits_NUM_BITS_5 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = 17'bxxxxxxxxxxxxxxxxx;
	rotated_data = _263;
end
always_comb begin // combinatorial offset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	offset_bits = 5'bxxxxx;
	offset_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 5'dx;
	_UIntToBits_value = offset;
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{17'bxxxxxxxxxxxxxxxxx, 17'bxxxxxxxxxxxxxxxxx, 17'bxxxxxxxxxxxxxxxxx, 17'bxxxxxxxxxxxxxxxxx, 17'bxxxxxxxxxxxxxxxxx, 17'bxxxxxxxxxxxxxxxxx};
	rotate_stages[0] = data;
	if(_4) rotate_stages[1][0] = _5;
	if(!_4) rotate_stages[1][0] = _6;
	if(_7) rotate_stages[1][1] = _8;
	if(!_7) rotate_stages[1][1] = _9;
	if(_10) rotate_stages[1][2] = _11;
	if(!_10) rotate_stages[1][2] = _12;
	if(_13) rotate_stages[1][3] = _14;
	if(!_13) rotate_stages[1][3] = _15;
	if(_16) rotate_stages[1][4] = _17;
	if(!_16) rotate_stages[1][4] = _18;
	if(_19) rotate_stages[1][5] = _20;
	if(!_19) rotate_stages[1][5] = _21;
	if(_22) rotate_stages[1][6] = _23;
	if(!_22) rotate_stages[1][6] = _24;
	if(_25) rotate_stages[1][7] = _26;
	if(!_25) rotate_stages[1][7] = _27;
	if(_28) rotate_stages[1][8] = _29;
	if(!_28) rotate_stages[1][8] = _30;
	if(_31) rotate_stages[1][9] = _32;
	if(!_31) rotate_stages[1][9] = _33;
	if(_34) rotate_stages[1][10] = _35;
	if(!_34) rotate_stages[1][10] = _36;
	if(_37) rotate_stages[1][11] = _38;
	if(!_37) rotate_stages[1][11] = _39;
	if(_40) rotate_stages[1][12] = _41;
	if(!_40) rotate_stages[1][12] = _42;
	if(_43) rotate_stages[1][13] = _44;
	if(!_43) rotate_stages[1][13] = _45;
	if(_46) rotate_stages[1][14] = _47;
	if(!_46) rotate_stages[1][14] = _48;
	if(_49) rotate_stages[1][15] = _50;
	if(!_49) rotate_stages[1][15] = _51;
	if(_52) rotate_stages[1][16] = _53;
	if(!_52) rotate_stages[1][16] = _54;
	if(_56) rotate_stages[2][0] = _57;
	if(!_56) rotate_stages[2][0] = _58;
	if(_59) rotate_stages[2][1] = _60;
	if(!_59) rotate_stages[2][1] = _61;
	if(_62) rotate_stages[2][2] = _63;
	if(!_62) rotate_stages[2][2] = _64;
	if(_65) rotate_stages[2][3] = _66;
	if(!_65) rotate_stages[2][3] = _67;
	if(_68) rotate_stages[2][4] = _69;
	if(!_68) rotate_stages[2][4] = _70;
	if(_71) rotate_stages[2][5] = _72;
	if(!_71) rotate_stages[2][5] = _73;
	if(_74) rotate_stages[2][6] = _75;
	if(!_74) rotate_stages[2][6] = _76;
	if(_77) rotate_stages[2][7] = _78;
	if(!_77) rotate_stages[2][7] = _79;
	if(_80) rotate_stages[2][8] = _81;
	if(!_80) rotate_stages[2][8] = _82;
	if(_83) rotate_stages[2][9] = _84;
	if(!_83) rotate_stages[2][9] = _85;
	if(_86) rotate_stages[2][10] = _87;
	if(!_86) rotate_stages[2][10] = _88;
	if(_89) rotate_stages[2][11] = _90;
	if(!_89) rotate_stages[2][11] = _91;
	if(_92) rotate_stages[2][12] = _93;
	if(!_92) rotate_stages[2][12] = _94;
	if(_95) rotate_stages[2][13] = _96;
	if(!_95) rotate_stages[2][13] = _97;
	if(_98) rotate_stages[2][14] = _99;
	if(!_98) rotate_stages[2][14] = _100;
	if(_101) rotate_stages[2][15] = _102;
	if(!_101) rotate_stages[2][15] = _103;
	if(_104) rotate_stages[2][16] = _105;
	if(!_104) rotate_stages[2][16] = _106;
	if(_108) rotate_stages[3][0] = _109;
	if(!_108) rotate_stages[3][0] = _110;
	if(_111) rotate_stages[3][1] = _112;
	if(!_111) rotate_stages[3][1] = _113;
	if(_114) rotate_stages[3][2] = _115;
	if(!_114) rotate_stages[3][2] = _116;
	if(_117) rotate_stages[3][3] = _118;
	if(!_117) rotate_stages[3][3] = _119;
	if(_120) rotate_stages[3][4] = _121;
	if(!_120) rotate_stages[3][4] = _122;
	if(_123) rotate_stages[3][5] = _124;
	if(!_123) rotate_stages[3][5] = _125;
	if(_126) rotate_stages[3][6] = _127;
	if(!_126) rotate_stages[3][6] = _128;
	if(_129) rotate_stages[3][7] = _130;
	if(!_129) rotate_stages[3][7] = _131;
	if(_132) rotate_stages[3][8] = _133;
	if(!_132) rotate_stages[3][8] = _134;
	if(_135) rotate_stages[3][9] = _136;
	if(!_135) rotate_stages[3][9] = _137;
	if(_138) rotate_stages[3][10] = _139;
	if(!_138) rotate_stages[3][10] = _140;
	if(_141) rotate_stages[3][11] = _142;
	if(!_141) rotate_stages[3][11] = _143;
	if(_144) rotate_stages[3][12] = _145;
	if(!_144) rotate_stages[3][12] = _146;
	if(_147) rotate_stages[3][13] = _148;
	if(!_147) rotate_stages[3][13] = _149;
	if(_150) rotate_stages[3][14] = _151;
	if(!_150) rotate_stages[3][14] = _152;
	if(_153) rotate_stages[3][15] = _154;
	if(!_153) rotate_stages[3][15] = _155;
	if(_156) rotate_stages[3][16] = _157;
	if(!_156) rotate_stages[3][16] = _158;
	if(_160) rotate_stages[4][0] = _161;
	if(!_160) rotate_stages[4][0] = _162;
	if(_163) rotate_stages[4][1] = _164;
	if(!_163) rotate_stages[4][1] = _165;
	if(_166) rotate_stages[4][2] = _167;
	if(!_166) rotate_stages[4][2] = _168;
	if(_169) rotate_stages[4][3] = _170;
	if(!_169) rotate_stages[4][3] = _171;
	if(_172) rotate_stages[4][4] = _173;
	if(!_172) rotate_stages[4][4] = _174;
	if(_175) rotate_stages[4][5] = _176;
	if(!_175) rotate_stages[4][5] = _177;
	if(_178) rotate_stages[4][6] = _179;
	if(!_178) rotate_stages[4][6] = _180;
	if(_181) rotate_stages[4][7] = _182;
	if(!_181) rotate_stages[4][7] = _183;
	if(_184) rotate_stages[4][8] = _185;
	if(!_184) rotate_stages[4][8] = _186;
	if(_187) rotate_stages[4][9] = _188;
	if(!_187) rotate_stages[4][9] = _189;
	if(_190) rotate_stages[4][10] = _191;
	if(!_190) rotate_stages[4][10] = _192;
	if(_193) rotate_stages[4][11] = _194;
	if(!_193) rotate_stages[4][11] = _195;
	if(_196) rotate_stages[4][12] = _197;
	if(!_196) rotate_stages[4][12] = _198;
	if(_199) rotate_stages[4][13] = _200;
	if(!_199) rotate_stages[4][13] = _201;
	if(_202) rotate_stages[4][14] = _203;
	if(!_202) rotate_stages[4][14] = _204;
	if(_205) rotate_stages[4][15] = _206;
	if(!_205) rotate_stages[4][15] = _207;
	if(_208) rotate_stages[4][16] = _209;
	if(!_208) rotate_stages[4][16] = _210;
	if(_212) rotate_stages[5][0] = _213;
	if(!_212) rotate_stages[5][0] = _214;
	if(_215) rotate_stages[5][1] = _216;
	if(!_215) rotate_stages[5][1] = _217;
	if(_218) rotate_stages[5][2] = _219;
	if(!_218) rotate_stages[5][2] = _220;
	if(_221) rotate_stages[5][3] = _222;
	if(!_221) rotate_stages[5][3] = _223;
	if(_224) rotate_stages[5][4] = _225;
	if(!_224) rotate_stages[5][4] = _226;
	if(_227) rotate_stages[5][5] = _228;
	if(!_227) rotate_stages[5][5] = _229;
	if(_230) rotate_stages[5][6] = _231;
	if(!_230) rotate_stages[5][6] = _232;
	if(_233) rotate_stages[5][7] = _234;
	if(!_233) rotate_stages[5][7] = _235;
	if(_236) rotate_stages[5][8] = _237;
	if(!_236) rotate_stages[5][8] = _238;
	if(_239) rotate_stages[5][9] = _240;
	if(!_239) rotate_stages[5][9] = _241;
	if(_242) rotate_stages[5][10] = _243;
	if(!_242) rotate_stages[5][10] = _244;
	if(_245) rotate_stages[5][11] = _246;
	if(!_245) rotate_stages[5][11] = _247;
	if(_248) rotate_stages[5][12] = _249;
	if(!_248) rotate_stages[5][12] = _250;
	if(_251) rotate_stages[5][13] = _252;
	if(!_251) rotate_stages[5][13] = _253;
	if(_254) rotate_stages[5][14] = _255;
	if(!_254) rotate_stages[5][14] = _256;
	if(_257) rotate_stages[5][15] = _258;
	if(!_257) rotate_stages[5][15] = _259;
	if(_260) rotate_stages[5][16] = _261;
	if(!_260) rotate_stages[5][16] = _262;
end
always_comb begin // combinatorial from
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from = 17'bxxxxxxxxxxxxxxxxx;
	from = _3;
end
always_comb begin // combinatorial from_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_2 = 17'bxxxxxxxxxxxxxxxxx;
	from_2 = _55;
end
always_comb begin // combinatorial from_3
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_3 = 17'bxxxxxxxxxxxxxxxxx;
	from_3 = _107;
end
always_comb begin // combinatorial from_4
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_4 = 17'bxxxxxxxxxxxxxxxxx;
	from_4 = _159;
end
always_comb begin // combinatorial from_5
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_5 = 17'bxxxxxxxxxxxxxxxxx;
	from_5 = _211;
end
endmodule

// RotateRight #(T: type bool #()[32], ARRAY_LEN: 17)
module RotateRight_T_type_bool_32_ARRAY_LEN_17(
	input clk,
	input wire[31:0] data[16:0],
	input wire[4:0] offset,
	output /*mux_wire*/ logic[31:0] rotated_data[16:0]
);

genvar _g0;
/*mux_wire*/ logic[4:0] offset_bits;
/*mux_wire*/ logic[4:0] _UIntToBits_value;
wire[4:0] _UIntToBits_bits;
/*mux_wire*/ logic[31:0] rotate_stages[5:0][16:0];
/*mux_wire*/ logic[31:0] from[16:0];
wire[31:0] _3[16:0];
generate
for(_g0 = 0; _g0 < 17; _g0 = _g0 + 1) begin
assign _3[_g0] = rotate_stages[0][_g0];
end
endgenerate
wire _4 = offset_bits[0];
wire[31:0] _5 = from[16];
wire[31:0] _6 = from[0];
wire _7 = offset_bits[0];
wire[31:0] _8 = from[0];
wire[31:0] _9 = from[1];
wire _10 = offset_bits[0];
wire[31:0] _11 = from[1];
wire[31:0] _12 = from[2];
wire _13 = offset_bits[0];
wire[31:0] _14 = from[2];
wire[31:0] _15 = from[3];
wire _16 = offset_bits[0];
wire[31:0] _17 = from[3];
wire[31:0] _18 = from[4];
wire _19 = offset_bits[0];
wire[31:0] _20 = from[4];
wire[31:0] _21 = from[5];
wire _22 = offset_bits[0];
wire[31:0] _23 = from[5];
wire[31:0] _24 = from[6];
wire _25 = offset_bits[0];
wire[31:0] _26 = from[6];
wire[31:0] _27 = from[7];
wire _28 = offset_bits[0];
wire[31:0] _29 = from[7];
wire[31:0] _30 = from[8];
wire _31 = offset_bits[0];
wire[31:0] _32 = from[8];
wire[31:0] _33 = from[9];
wire _34 = offset_bits[0];
wire[31:0] _35 = from[9];
wire[31:0] _36 = from[10];
wire _37 = offset_bits[0];
wire[31:0] _38 = from[10];
wire[31:0] _39 = from[11];
wire _40 = offset_bits[0];
wire[31:0] _41 = from[11];
wire[31:0] _42 = from[12];
wire _43 = offset_bits[0];
wire[31:0] _44 = from[12];
wire[31:0] _45 = from[13];
wire _46 = offset_bits[0];
wire[31:0] _47 = from[13];
wire[31:0] _48 = from[14];
wire _49 = offset_bits[0];
wire[31:0] _50 = from[14];
wire[31:0] _51 = from[15];
wire _52 = offset_bits[0];
wire[31:0] _53 = from[15];
wire[31:0] _54 = from[16];
/*mux_wire*/ logic[31:0] from_2[16:0];
wire[31:0] _55[16:0];
generate
for(_g0 = 0; _g0 < 17; _g0 = _g0 + 1) begin
assign _55[_g0] = rotate_stages[1][_g0];
end
endgenerate
wire _56 = offset_bits[1];
wire[31:0] _57 = from_2[15];
wire[31:0] _58 = from_2[0];
wire _59 = offset_bits[1];
wire[31:0] _60 = from_2[16];
wire[31:0] _61 = from_2[1];
wire _62 = offset_bits[1];
wire[31:0] _63 = from_2[0];
wire[31:0] _64 = from_2[2];
wire _65 = offset_bits[1];
wire[31:0] _66 = from_2[1];
wire[31:0] _67 = from_2[3];
wire _68 = offset_bits[1];
wire[31:0] _69 = from_2[2];
wire[31:0] _70 = from_2[4];
wire _71 = offset_bits[1];
wire[31:0] _72 = from_2[3];
wire[31:0] _73 = from_2[5];
wire _74 = offset_bits[1];
wire[31:0] _75 = from_2[4];
wire[31:0] _76 = from_2[6];
wire _77 = offset_bits[1];
wire[31:0] _78 = from_2[5];
wire[31:0] _79 = from_2[7];
wire _80 = offset_bits[1];
wire[31:0] _81 = from_2[6];
wire[31:0] _82 = from_2[8];
wire _83 = offset_bits[1];
wire[31:0] _84 = from_2[7];
wire[31:0] _85 = from_2[9];
wire _86 = offset_bits[1];
wire[31:0] _87 = from_2[8];
wire[31:0] _88 = from_2[10];
wire _89 = offset_bits[1];
wire[31:0] _90 = from_2[9];
wire[31:0] _91 = from_2[11];
wire _92 = offset_bits[1];
wire[31:0] _93 = from_2[10];
wire[31:0] _94 = from_2[12];
wire _95 = offset_bits[1];
wire[31:0] _96 = from_2[11];
wire[31:0] _97 = from_2[13];
wire _98 = offset_bits[1];
wire[31:0] _99 = from_2[12];
wire[31:0] _100 = from_2[14];
wire _101 = offset_bits[1];
wire[31:0] _102 = from_2[13];
wire[31:0] _103 = from_2[15];
wire _104 = offset_bits[1];
wire[31:0] _105 = from_2[14];
wire[31:0] _106 = from_2[16];
/*mux_wire*/ logic[31:0] from_3[16:0];
wire[31:0] _107[16:0];
generate
for(_g0 = 0; _g0 < 17; _g0 = _g0 + 1) begin
assign _107[_g0] = rotate_stages[2][_g0];
end
endgenerate
wire _108 = offset_bits[2];
wire[31:0] _109 = from_3[13];
wire[31:0] _110 = from_3[0];
wire _111 = offset_bits[2];
wire[31:0] _112 = from_3[14];
wire[31:0] _113 = from_3[1];
wire _114 = offset_bits[2];
wire[31:0] _115 = from_3[15];
wire[31:0] _116 = from_3[2];
wire _117 = offset_bits[2];
wire[31:0] _118 = from_3[16];
wire[31:0] _119 = from_3[3];
wire _120 = offset_bits[2];
wire[31:0] _121 = from_3[0];
wire[31:0] _122 = from_3[4];
wire _123 = offset_bits[2];
wire[31:0] _124 = from_3[1];
wire[31:0] _125 = from_3[5];
wire _126 = offset_bits[2];
wire[31:0] _127 = from_3[2];
wire[31:0] _128 = from_3[6];
wire _129 = offset_bits[2];
wire[31:0] _130 = from_3[3];
wire[31:0] _131 = from_3[7];
wire _132 = offset_bits[2];
wire[31:0] _133 = from_3[4];
wire[31:0] _134 = from_3[8];
wire _135 = offset_bits[2];
wire[31:0] _136 = from_3[5];
wire[31:0] _137 = from_3[9];
wire _138 = offset_bits[2];
wire[31:0] _139 = from_3[6];
wire[31:0] _140 = from_3[10];
wire _141 = offset_bits[2];
wire[31:0] _142 = from_3[7];
wire[31:0] _143 = from_3[11];
wire _144 = offset_bits[2];
wire[31:0] _145 = from_3[8];
wire[31:0] _146 = from_3[12];
wire _147 = offset_bits[2];
wire[31:0] _148 = from_3[9];
wire[31:0] _149 = from_3[13];
wire _150 = offset_bits[2];
wire[31:0] _151 = from_3[10];
wire[31:0] _152 = from_3[14];
wire _153 = offset_bits[2];
wire[31:0] _154 = from_3[11];
wire[31:0] _155 = from_3[15];
wire _156 = offset_bits[2];
wire[31:0] _157 = from_3[12];
wire[31:0] _158 = from_3[16];
/*mux_wire*/ logic[31:0] from_4[16:0];
wire[31:0] _159[16:0];
generate
for(_g0 = 0; _g0 < 17; _g0 = _g0 + 1) begin
assign _159[_g0] = rotate_stages[3][_g0];
end
endgenerate
wire _160 = offset_bits[3];
wire[31:0] _161 = from_4[9];
wire[31:0] _162 = from_4[0];
wire _163 = offset_bits[3];
wire[31:0] _164 = from_4[10];
wire[31:0] _165 = from_4[1];
wire _166 = offset_bits[3];
wire[31:0] _167 = from_4[11];
wire[31:0] _168 = from_4[2];
wire _169 = offset_bits[3];
wire[31:0] _170 = from_4[12];
wire[31:0] _171 = from_4[3];
wire _172 = offset_bits[3];
wire[31:0] _173 = from_4[13];
wire[31:0] _174 = from_4[4];
wire _175 = offset_bits[3];
wire[31:0] _176 = from_4[14];
wire[31:0] _177 = from_4[5];
wire _178 = offset_bits[3];
wire[31:0] _179 = from_4[15];
wire[31:0] _180 = from_4[6];
wire _181 = offset_bits[3];
wire[31:0] _182 = from_4[16];
wire[31:0] _183 = from_4[7];
wire _184 = offset_bits[3];
wire[31:0] _185 = from_4[0];
wire[31:0] _186 = from_4[8];
wire _187 = offset_bits[3];
wire[31:0] _188 = from_4[1];
wire[31:0] _189 = from_4[9];
wire _190 = offset_bits[3];
wire[31:0] _191 = from_4[2];
wire[31:0] _192 = from_4[10];
wire _193 = offset_bits[3];
wire[31:0] _194 = from_4[3];
wire[31:0] _195 = from_4[11];
wire _196 = offset_bits[3];
wire[31:0] _197 = from_4[4];
wire[31:0] _198 = from_4[12];
wire _199 = offset_bits[3];
wire[31:0] _200 = from_4[5];
wire[31:0] _201 = from_4[13];
wire _202 = offset_bits[3];
wire[31:0] _203 = from_4[6];
wire[31:0] _204 = from_4[14];
wire _205 = offset_bits[3];
wire[31:0] _206 = from_4[7];
wire[31:0] _207 = from_4[15];
wire _208 = offset_bits[3];
wire[31:0] _209 = from_4[8];
wire[31:0] _210 = from_4[16];
/*mux_wire*/ logic[31:0] from_5[16:0];
wire[31:0] _211[16:0];
generate
for(_g0 = 0; _g0 < 17; _g0 = _g0 + 1) begin
assign _211[_g0] = rotate_stages[4][_g0];
end
endgenerate
wire _212 = offset_bits[4];
wire[31:0] _213 = from_5[1];
wire[31:0] _214 = from_5[0];
wire _215 = offset_bits[4];
wire[31:0] _216 = from_5[2];
wire[31:0] _217 = from_5[1];
wire _218 = offset_bits[4];
wire[31:0] _219 = from_5[3];
wire[31:0] _220 = from_5[2];
wire _221 = offset_bits[4];
wire[31:0] _222 = from_5[4];
wire[31:0] _223 = from_5[3];
wire _224 = offset_bits[4];
wire[31:0] _225 = from_5[5];
wire[31:0] _226 = from_5[4];
wire _227 = offset_bits[4];
wire[31:0] _228 = from_5[6];
wire[31:0] _229 = from_5[5];
wire _230 = offset_bits[4];
wire[31:0] _231 = from_5[7];
wire[31:0] _232 = from_5[6];
wire _233 = offset_bits[4];
wire[31:0] _234 = from_5[8];
wire[31:0] _235 = from_5[7];
wire _236 = offset_bits[4];
wire[31:0] _237 = from_5[9];
wire[31:0] _238 = from_5[8];
wire _239 = offset_bits[4];
wire[31:0] _240 = from_5[10];
wire[31:0] _241 = from_5[9];
wire _242 = offset_bits[4];
wire[31:0] _243 = from_5[11];
wire[31:0] _244 = from_5[10];
wire _245 = offset_bits[4];
wire[31:0] _246 = from_5[12];
wire[31:0] _247 = from_5[11];
wire _248 = offset_bits[4];
wire[31:0] _249 = from_5[13];
wire[31:0] _250 = from_5[12];
wire _251 = offset_bits[4];
wire[31:0] _252 = from_5[14];
wire[31:0] _253 = from_5[13];
wire _254 = offset_bits[4];
wire[31:0] _255 = from_5[15];
wire[31:0] _256 = from_5[14];
wire _257 = offset_bits[4];
wire[31:0] _258 = from_5[16];
wire[31:0] _259 = from_5[15];
wire _260 = offset_bits[4];
wire[31:0] _261 = from_5[0];
wire[31:0] _262 = from_5[16];
wire[31:0] _263[16:0];
generate
for(_g0 = 0; _g0 < 17; _g0 = _g0 + 1) begin
assign _263[_g0] = rotate_stages[5][_g0];
end
endgenerate
UIntToBits_NUM_BITS_5 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
always_comb begin // combinatorial rotated_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotated_data = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 17; _v0 = _v0 + 1) begin
rotated_data[_v0] = _263[_v0];
end
end
always_comb begin // combinatorial offset_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	offset_bits = 5'bxxxxx;
	offset_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 5'dx;
	_UIntToBits_value = offset;
end
always_comb begin // combinatorial rotate_stages
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rotate_stages = '{'{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}, '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx}};
	for(int _v0 = 0; _v0 < 17; _v0 = _v0 + 1) begin
rotate_stages[0][_v0] = data[_v0];
end
	if(_4) rotate_stages[1][0] = _5;
	if(!_4) rotate_stages[1][0] = _6;
	if(_7) rotate_stages[1][1] = _8;
	if(!_7) rotate_stages[1][1] = _9;
	if(_10) rotate_stages[1][2] = _11;
	if(!_10) rotate_stages[1][2] = _12;
	if(_13) rotate_stages[1][3] = _14;
	if(!_13) rotate_stages[1][3] = _15;
	if(_16) rotate_stages[1][4] = _17;
	if(!_16) rotate_stages[1][4] = _18;
	if(_19) rotate_stages[1][5] = _20;
	if(!_19) rotate_stages[1][5] = _21;
	if(_22) rotate_stages[1][6] = _23;
	if(!_22) rotate_stages[1][6] = _24;
	if(_25) rotate_stages[1][7] = _26;
	if(!_25) rotate_stages[1][7] = _27;
	if(_28) rotate_stages[1][8] = _29;
	if(!_28) rotate_stages[1][8] = _30;
	if(_31) rotate_stages[1][9] = _32;
	if(!_31) rotate_stages[1][9] = _33;
	if(_34) rotate_stages[1][10] = _35;
	if(!_34) rotate_stages[1][10] = _36;
	if(_37) rotate_stages[1][11] = _38;
	if(!_37) rotate_stages[1][11] = _39;
	if(_40) rotate_stages[1][12] = _41;
	if(!_40) rotate_stages[1][12] = _42;
	if(_43) rotate_stages[1][13] = _44;
	if(!_43) rotate_stages[1][13] = _45;
	if(_46) rotate_stages[1][14] = _47;
	if(!_46) rotate_stages[1][14] = _48;
	if(_49) rotate_stages[1][15] = _50;
	if(!_49) rotate_stages[1][15] = _51;
	if(_52) rotate_stages[1][16] = _53;
	if(!_52) rotate_stages[1][16] = _54;
	if(_56) rotate_stages[2][0] = _57;
	if(!_56) rotate_stages[2][0] = _58;
	if(_59) rotate_stages[2][1] = _60;
	if(!_59) rotate_stages[2][1] = _61;
	if(_62) rotate_stages[2][2] = _63;
	if(!_62) rotate_stages[2][2] = _64;
	if(_65) rotate_stages[2][3] = _66;
	if(!_65) rotate_stages[2][3] = _67;
	if(_68) rotate_stages[2][4] = _69;
	if(!_68) rotate_stages[2][4] = _70;
	if(_71) rotate_stages[2][5] = _72;
	if(!_71) rotate_stages[2][5] = _73;
	if(_74) rotate_stages[2][6] = _75;
	if(!_74) rotate_stages[2][6] = _76;
	if(_77) rotate_stages[2][7] = _78;
	if(!_77) rotate_stages[2][7] = _79;
	if(_80) rotate_stages[2][8] = _81;
	if(!_80) rotate_stages[2][8] = _82;
	if(_83) rotate_stages[2][9] = _84;
	if(!_83) rotate_stages[2][9] = _85;
	if(_86) rotate_stages[2][10] = _87;
	if(!_86) rotate_stages[2][10] = _88;
	if(_89) rotate_stages[2][11] = _90;
	if(!_89) rotate_stages[2][11] = _91;
	if(_92) rotate_stages[2][12] = _93;
	if(!_92) rotate_stages[2][12] = _94;
	if(_95) rotate_stages[2][13] = _96;
	if(!_95) rotate_stages[2][13] = _97;
	if(_98) rotate_stages[2][14] = _99;
	if(!_98) rotate_stages[2][14] = _100;
	if(_101) rotate_stages[2][15] = _102;
	if(!_101) rotate_stages[2][15] = _103;
	if(_104) rotate_stages[2][16] = _105;
	if(!_104) rotate_stages[2][16] = _106;
	if(_108) rotate_stages[3][0] = _109;
	if(!_108) rotate_stages[3][0] = _110;
	if(_111) rotate_stages[3][1] = _112;
	if(!_111) rotate_stages[3][1] = _113;
	if(_114) rotate_stages[3][2] = _115;
	if(!_114) rotate_stages[3][2] = _116;
	if(_117) rotate_stages[3][3] = _118;
	if(!_117) rotate_stages[3][3] = _119;
	if(_120) rotate_stages[3][4] = _121;
	if(!_120) rotate_stages[3][4] = _122;
	if(_123) rotate_stages[3][5] = _124;
	if(!_123) rotate_stages[3][5] = _125;
	if(_126) rotate_stages[3][6] = _127;
	if(!_126) rotate_stages[3][6] = _128;
	if(_129) rotate_stages[3][7] = _130;
	if(!_129) rotate_stages[3][7] = _131;
	if(_132) rotate_stages[3][8] = _133;
	if(!_132) rotate_stages[3][8] = _134;
	if(_135) rotate_stages[3][9] = _136;
	if(!_135) rotate_stages[3][9] = _137;
	if(_138) rotate_stages[3][10] = _139;
	if(!_138) rotate_stages[3][10] = _140;
	if(_141) rotate_stages[3][11] = _142;
	if(!_141) rotate_stages[3][11] = _143;
	if(_144) rotate_stages[3][12] = _145;
	if(!_144) rotate_stages[3][12] = _146;
	if(_147) rotate_stages[3][13] = _148;
	if(!_147) rotate_stages[3][13] = _149;
	if(_150) rotate_stages[3][14] = _151;
	if(!_150) rotate_stages[3][14] = _152;
	if(_153) rotate_stages[3][15] = _154;
	if(!_153) rotate_stages[3][15] = _155;
	if(_156) rotate_stages[3][16] = _157;
	if(!_156) rotate_stages[3][16] = _158;
	if(_160) rotate_stages[4][0] = _161;
	if(!_160) rotate_stages[4][0] = _162;
	if(_163) rotate_stages[4][1] = _164;
	if(!_163) rotate_stages[4][1] = _165;
	if(_166) rotate_stages[4][2] = _167;
	if(!_166) rotate_stages[4][2] = _168;
	if(_169) rotate_stages[4][3] = _170;
	if(!_169) rotate_stages[4][3] = _171;
	if(_172) rotate_stages[4][4] = _173;
	if(!_172) rotate_stages[4][4] = _174;
	if(_175) rotate_stages[4][5] = _176;
	if(!_175) rotate_stages[4][5] = _177;
	if(_178) rotate_stages[4][6] = _179;
	if(!_178) rotate_stages[4][6] = _180;
	if(_181) rotate_stages[4][7] = _182;
	if(!_181) rotate_stages[4][7] = _183;
	if(_184) rotate_stages[4][8] = _185;
	if(!_184) rotate_stages[4][8] = _186;
	if(_187) rotate_stages[4][9] = _188;
	if(!_187) rotate_stages[4][9] = _189;
	if(_190) rotate_stages[4][10] = _191;
	if(!_190) rotate_stages[4][10] = _192;
	if(_193) rotate_stages[4][11] = _194;
	if(!_193) rotate_stages[4][11] = _195;
	if(_196) rotate_stages[4][12] = _197;
	if(!_196) rotate_stages[4][12] = _198;
	if(_199) rotate_stages[4][13] = _200;
	if(!_199) rotate_stages[4][13] = _201;
	if(_202) rotate_stages[4][14] = _203;
	if(!_202) rotate_stages[4][14] = _204;
	if(_205) rotate_stages[4][15] = _206;
	if(!_205) rotate_stages[4][15] = _207;
	if(_208) rotate_stages[4][16] = _209;
	if(!_208) rotate_stages[4][16] = _210;
	if(_212) rotate_stages[5][0] = _213;
	if(!_212) rotate_stages[5][0] = _214;
	if(_215) rotate_stages[5][1] = _216;
	if(!_215) rotate_stages[5][1] = _217;
	if(_218) rotate_stages[5][2] = _219;
	if(!_218) rotate_stages[5][2] = _220;
	if(_221) rotate_stages[5][3] = _222;
	if(!_221) rotate_stages[5][3] = _223;
	if(_224) rotate_stages[5][4] = _225;
	if(!_224) rotate_stages[5][4] = _226;
	if(_227) rotate_stages[5][5] = _228;
	if(!_227) rotate_stages[5][5] = _229;
	if(_230) rotate_stages[5][6] = _231;
	if(!_230) rotate_stages[5][6] = _232;
	if(_233) rotate_stages[5][7] = _234;
	if(!_233) rotate_stages[5][7] = _235;
	if(_236) rotate_stages[5][8] = _237;
	if(!_236) rotate_stages[5][8] = _238;
	if(_239) rotate_stages[5][9] = _240;
	if(!_239) rotate_stages[5][9] = _241;
	if(_242) rotate_stages[5][10] = _243;
	if(!_242) rotate_stages[5][10] = _244;
	if(_245) rotate_stages[5][11] = _246;
	if(!_245) rotate_stages[5][11] = _247;
	if(_248) rotate_stages[5][12] = _249;
	if(!_248) rotate_stages[5][12] = _250;
	if(_251) rotate_stages[5][13] = _252;
	if(!_251) rotate_stages[5][13] = _253;
	if(_254) rotate_stages[5][14] = _255;
	if(!_254) rotate_stages[5][14] = _256;
	if(_257) rotate_stages[5][15] = _258;
	if(!_257) rotate_stages[5][15] = _259;
	if(_260) rotate_stages[5][16] = _261;
	if(!_260) rotate_stages[5][16] = _262;
end
always_comb begin // combinatorial from
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 17; _v0 = _v0 + 1) begin
from[_v0] = _3[_v0];
end
end
always_comb begin // combinatorial from_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_2 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 17; _v0 = _v0 + 1) begin
from_2[_v0] = _55[_v0];
end
end
always_comb begin // combinatorial from_3
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_3 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 17; _v0 = _v0 + 1) begin
from_3[_v0] = _107[_v0];
end
end
always_comb begin // combinatorial from_4
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_4 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 17; _v0 = _v0 + 1) begin
from_4[_v0] = _159[_v0];
end
end
always_comb begin // combinatorial from_5
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	from_5 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 17; _v0 = _v0 + 1) begin
from_5[_v0] = _211[_v0];
end
end
endmodule

// UIntToBits #(NUM_BITS: 5)
module UIntToBits_NUM_BITS_5(
	input clk,
	input wire[4:0] value,
	output /*mux_wire*/ logic[4:0] bits
);

	assign bits = value;
endmodule

// axi_array_burst_reader #(AXI_WIDTH: 512, ADDR_ALIGN: 4, COUNT_TO: 1114112, ATO: 18446744073709551616)
module axi_array_burst_reader_AXI_WIDTH_512_ADDR_ALIGN_4_COUNT_TO_1114112_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*state*/ logic arvalid,
	input wire arready,
	output /*state*/ logic[63:0] araddr,
	output /*state*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[511:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic element_packet_valid,
	output /*mux_wire*/ logic[31:0] elements[15:0],
	output /*mux_wire*/ logic[3:0] chunk_offset,
	output /*mux_wire*/ logic[4:0] chunk_length,
	output /*mux_wire*/ logic last,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[20:0] count
);

/*latency*/ logic _arvalid_D1; always_ff @(posedge aclk) begin _arvalid_D1 <= arvalid; end
/*latency*/ logic _request_new_burst_D1; always_ff @(posedge aclk) begin _request_new_burst_D1 <= request_new_burst; end
genvar _g0;
localparam[1:0] _1 = 2'b01;
localparam[2:0] _2 = 3'b000;
localparam[3:0] _3 = 4'b0010;
/*mux_wire*/ logic[1:0] _rresp;
/*mux_wire*/ logic _rlast;
/*state*/ logic[11:0] num_in_flight;
/*state*/ logic last_burst_in_flight;
/*mux_wire*/ logic[63:0] next_araddr;
/*latency*/ logic[63:0] _next_araddr_D0; always_ff @(posedge aclk) begin _next_araddr_D0 <= next_araddr; end
wire[57:0] _cur_start_chunk_addr_old;
/*mux_wire*/ logic[57:0] _BitwiseIntConcat_upper;
/*mux_wire*/ logic[5:0] _BitwiseIntConcat_lower;
wire[63:0] _BitwiseIntConcat_v;
/*mux_wire*/ logic[5:0] next_arlen;
/*mux_wire*/ logic next_last_burst_in_flight;
/*latency*/ logic _next_last_burst_in_flight_D0; always_ff @(posedge aclk) begin _next_last_burst_in_flight_D0 <= next_last_burst_in_flight; end
/*mux_wire*/ logic[51:0] cur_burst_addr;
/*mux_wire*/ logic[5:0] cur_align;
/*mux_wire*/ logic[57:0] _BitwiseIntSplit_v;
wire[51:0] _BitwiseIntSplit_upper;
wire[5:0] _BitwiseIntSplit_lower;
/*mux_wire*/ logic chunks_are_left;
/*latency*/ logic _chunks_are_left_D0; always_ff @(posedge aclk) begin _chunks_are_left_D0 <= chunks_are_left; end
wire[16:0] _num_chunks_left_old;
/*latency*/ logic[16:0] __num_chunks_left_old_N1; always_ff @(posedge aclk) begin __num_chunks_left_old_N1 <= _num_chunks_left_old; end
/*latency*/ logic[16:0] __num_chunks_left_old_D0; always_ff @(posedge aclk) begin __num_chunks_left_old_D0 <= __num_chunks_left_old_N1; end
wire _14;
assign _14 = _num_chunks_left_old > 1'd0;
/*latency*/ logic __14_N1; always_ff @(posedge aclk) begin __14_N1 <= _14; end
/*mux_wire*/ logic[5:0] max_chunks_in_this_burst;
/*latency*/ logic[5:0] _max_chunks_in_this_burst_D0; always_ff @(posedge aclk) begin _max_chunks_in_this_burst_D0 <= max_chunks_in_this_burst; end
wire[5:0] _18;
assign _18 = 6'd63 - cur_align;
wire[6:0] _22;
assign _22 = max_chunks_in_this_burst + 1'd1;
wire _23;
assign _23 = __num_chunks_left_old_N1 <= _22;
/*latency*/ logic __23_D0; always_ff @(posedge aclk) begin __23_D0 <= _23; end
/*mux_wire*/ logic[16:0] _IntNarrow_in;
wire[6:0] _IntNarrow_out;
wire[5:0] _26;
assign _26 = _IntNarrow_out - 1'd1;
/*latency*/ logic[5:0] __26_D0; always_ff @(posedge aclk) begin __26_D0 <= _26; end
/*mux_wire*/ logic may_next_arvalid;
/*latency*/ logic _may_next_arvalid_D1; always_ff @(posedge aclk) begin _may_next_arvalid_D1 <= may_next_arvalid; end
wire _num_chunks_left_may_update;
wire _30;
assign _30 = _chunks_are_left_D0 & _num_chunks_left_may_update;
wire _cur_start_chunk_addr_may_update;
wire _32;
assign _32 = _30 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
wire _34;
assign _34 = _32 & _LatencyOffset_out;
wire signed[11:0] _37;
assign _37 = max_in_flight - 7'd64;
wire _38;
assign _38 = $signed({1'b0, num_in_flight}) <= _37;
wire _39;
assign _39 = _34 & _38;
/*mux_wire*/ logic[52:0] next_burst_addr;
wire[52:0] _45;
assign _45 = cur_burst_addr + 1'd1;
/*latency*/ logic[52:0] __45_D0; always_ff @(posedge aclk) begin __45_D0 <= _45; end
/*latency*/ logic[52:0] __45_D1; always_ff @(posedge aclk) begin __45_D1 <= __45_D0; end
/*mux_wire*/ logic[52:0] _BitwiseIntConcat_2_upper;
/*mux_wire*/ logic[5:0] _BitwiseIntConcat_2_lower;
wire[58:0] _BitwiseIntConcat_2_v;
/*mux_wire*/ logic[58:0] _IntNarrow_2_in;
wire[57:0] _IntNarrow_2_out;
/*mux_wire*/ logic _cur_start_chunk_addr_update;
/*mux_wire*/ logic[57:0] _cur_start_chunk_addr_new;
/*mux_wire*/ logic[16:0] next_num_chunks_left;
wire[6:0] _53;
assign _53 = next_arlen + 1'd1;
wire signed[17:0] _54;
assign _54 = __num_chunks_left_old_D0 - _53;
/*mux_wire*/ logic signed[17:0] _IntNarrow_3_in;
wire[16:0] _IntNarrow_3_out;
/*mux_wire*/ logic _num_chunks_left_update;
/*mux_wire*/ logic[16:0] _num_chunks_left_new;
/*mux_wire*/ logic _BoolToInt_i;
wire[0:0] _BoolToInt_o;
wire signed[12:0] _64;
assign _64 = num_in_flight - _BoolToInt_o;
wire _66;
assign _66 = !arvalid;
wire _68;
assign _68 = _66 & may_next_arvalid;
wire[6:0] _71;
assign _71 = next_arlen + 1'd1;
/*mux_wire*/ logic _Ternary_cond;
/*mux_wire*/ logic[6:0] _Ternary_a;
/*mux_wire*/ logic[6:0] _Ternary_b;
wire[6:0] _Ternary_o;
wire signed[12:0] _73;
assign _73 = _64 + $signed({1'b0, _Ternary_o});
/*mux_wire*/ logic signed[12:0] _IntNarrow_4_in;
wire[11:0] _IntNarrow_4_out;
/*state*/ logic[4:0] final_chunk_align;
/*state*/ logic[3:0] cur_chunk_align;
/*mux_wire*/ logic[31:0] elements_2[15:0];
wire[31:0] _75;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _75[_g0] = rdata[_g0];
end
endgenerate
wire[31:0] _76;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _76[_g0] = rdata[32 + _g0];
end
endgenerate
wire[31:0] _77;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _77[_g0] = rdata[64 + _g0];
end
endgenerate
wire[31:0] _78;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _78[_g0] = rdata[96 + _g0];
end
endgenerate
wire[31:0] _79;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _79[_g0] = rdata[128 + _g0];
end
endgenerate
wire[31:0] _80;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _80[_g0] = rdata[160 + _g0];
end
endgenerate
wire[31:0] _81;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _81[_g0] = rdata[192 + _g0];
end
endgenerate
wire[31:0] _82;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _82[_g0] = rdata[224 + _g0];
end
endgenerate
wire[31:0] _83;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _83[_g0] = rdata[256 + _g0];
end
endgenerate
wire[31:0] _84;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _84[_g0] = rdata[288 + _g0];
end
endgenerate
wire[31:0] _85;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _85[_g0] = rdata[320 + _g0];
end
endgenerate
wire[31:0] _86;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _86[_g0] = rdata[352 + _g0];
end
endgenerate
wire[31:0] _87;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _87[_g0] = rdata[384 + _g0];
end
endgenerate
wire[31:0] _88;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _88[_g0] = rdata[416 + _g0];
end
endgenerate
wire[31:0] _89;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _89[_g0] = rdata[448 + _g0];
end
endgenerate
wire[31:0] _90;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _90[_g0] = rdata[480 + _g0];
end
endgenerate
/*mux_wire*/ logic[4:0] num_chunk_elements;
/*mux_wire*/ logic is_last;
wire _93;
assign _93 = num_in_flight == 1'd1;
wire _95;
assign _95 = _93 & last_burst_in_flight;
wire signed[5:0] _99;
assign _99 = final_chunk_align - cur_chunk_align;
/*mux_wire*/ logic signed[5:0] _IntNarrow_5_in;
wire[4:0] _IntNarrow_5_out;
wire[4:0] _101;
assign _101 = 5'd16 - cur_chunk_align;
wire _109;
assign _109 = !chunks_are_left;
/*latency*/ logic __109_D0; always_ff @(posedge aclk) begin __109_D0 <= _109; end
wire _111;
assign _111 = __109_D0 & _num_chunks_left_may_update;
wire _113;
assign _113 = _111 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic[57:0] chunk_addr;
/*latency*/ logic[57:0] _chunk_addr_D1; always_ff @(posedge aclk) begin _chunk_addr_D1 <= chunk_addr; end
/*mux_wire*/ logic[3:0] element_in_chunk_align;
wire[61:0] _115;
assign _115 = start_addr / 3'd4;
/*mux_wire*/ logic[61:0] _BitwiseIntSplit_2_v;
wire[57:0] _BitwiseIntSplit_2_upper;
wire[3:0] _BitwiseIntSplit_2_lower;
/*mux_wire*/ logic[16:0] chunk_count_bits;
/*mux_wire*/ logic[3:0] final_alignment;
wire[20:0] _118;
assign _118 = count + element_in_chunk_align;
/*mux_wire*/ logic[20:0] _BitwiseIntSplit_3_v;
wire[16:0] _BitwiseIntSplit_3_upper;
wire[3:0] _BitwiseIntSplit_3_lower;
/*mux_wire*/ logic[16:0] num_chunks;
/*mux_wire*/ logic is_no_chunks;
wire _121;
assign _121 = chunk_count_bits == 1'd0;
wire _127;
assign _127 = final_alignment != 1'd0;
/*mux_wire*/ logic _BoolToInt_2_i;
wire[0:0] _BoolToInt_2_o;
wire[16:0] _128;
assign _128 = chunk_count_bits + _BoolToInt_2_o;
wire _134;
assign _134 = !is_no_chunks;
wire _137;
assign _137 = final_alignment == 1'd0;
wire _138;
assign _138 = _134 & _137;
/*mux_wire*/ logic _BoolToInt_3_i;
wire[0:0] _BoolToInt_3_o;
/*mux_wire*/ logic[0:0] _BitwiseIntConcat_3_upper;
/*mux_wire*/ logic[3:0] _BitwiseIntConcat_3_lower;
wire[4:0] _BitwiseIntConcat_3_v;
wire _142;
assign _142 = !aresetn;
/*mux_wire*/ logic _cur_start_chunk_addr_rst;
wire _144;
assign _144 = !aresetn;
/*mux_wire*/ logic _num_chunks_left_rst;
wire _146;
assign _146 = !aresetn;
SlowState_T_type_int_FROM_0_TO_288230376151711744_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1 cur_start_chunk_addr(
	.clk(aclk),
	.rst(_cur_start_chunk_addr_rst),
	.old(_cur_start_chunk_addr_old),
	.may_update(_cur_start_chunk_addr_may_update),
	.update(_cur_start_chunk_addr_update),
	.new_1(_cur_start_chunk_addr_new)
);
SlowState_T_type_int_FROM_0_TO_69635_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0 num_chunks_left(
	.clk(aclk),
	.rst(_num_chunks_left_rst),
	.old(_num_chunks_left_old),
	.may_update(_num_chunks_left_may_update),
	.update(_num_chunks_left_update),
	.new_1(_num_chunks_left_new)
);
BitwiseIntConcat_UPPER_TO_288230376151711744_LOWER_BITS_6 BitwiseIntConcat(
	.clk(aclk),
	.upper(_BitwiseIntConcat_upper),
	.lower(_BitwiseIntConcat_lower),
	.v(_BitwiseIntConcat_v)
);
BitwiseIntSplit_TO_288230376151711744_LOWER_BITS_6 BitwiseIntSplit(
	.clk(aclk),
	.v(_BitwiseIntSplit_v),
	.upper(_BitwiseIntSplit_upper),
	.lower(_BitwiseIntSplit_lower)
);
IntNarrow_FROM_I_0_TO_I_69635_FROM_1_TO_65 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
LatencyOffset_T_type_bool_OFFSET_192 LatencyOffset(
	.clk(aclk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
BitwiseIntConcat_UPPER_TO_4503599627370497_LOWER_BITS_6 BitwiseIntConcat_2(
	.clk(aclk),
	.upper(_BitwiseIntConcat_2_upper),
	.lower(_BitwiseIntConcat_2_lower),
	.v(_BitwiseIntConcat_2_v)
);
IntNarrow_FROM_I_0_TO_I_288230376151711808_FROM_0_TO_288230376151711744 IntNarrow_2(
	.clk(aclk),
	.in(_IntNarrow_2_in),
	.out(_IntNarrow_2_out)
);
IntNarrow_FROM_I_64_TO_I_69634_FROM_0_TO_69635 IntNarrow_3(
	.clk(aclk),
	.in(_IntNarrow_3_in),
	.out(_IntNarrow_3_out)
);
BoolToInt BoolToInt(
	.clk(aclk),
	.i(_BoolToInt_i),
	.o(_BoolToInt_o)
);
Ternary_T_type_int_FROM_0_TO_65 Ternary(
	.clk(aclk),
	.cond(_Ternary_cond),
	.a(_Ternary_a),
	.b(_Ternary_b),
	.o(_Ternary_o)
);
IntNarrow_FROM_I_1_TO_I_3256_FROM_0_TO_3192 IntNarrow_4(
	.clk(aclk),
	.in(_IntNarrow_4_in),
	.out(_IntNarrow_4_out)
);
IntNarrow_FROM_I_15_TO_I_32_FROM_0_TO_17 IntNarrow_5(
	.clk(aclk),
	.in(_IntNarrow_5_in),
	.out(_IntNarrow_5_out)
);
BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_4 BitwiseIntSplit_2(
	.clk(aclk),
	.v(_BitwiseIntSplit_2_v),
	.upper(_BitwiseIntSplit_2_upper),
	.lower(_BitwiseIntSplit_2_lower)
);
BitwiseIntSplit_TO_1114127_LOWER_BITS_4 BitwiseIntSplit_3(
	.clk(aclk),
	.v(_BitwiseIntSplit_3_v),
	.upper(_BitwiseIntSplit_3_upper),
	.lower(_BitwiseIntSplit_3_lower)
);
BoolToInt BoolToInt_2(
	.clk(aclk),
	.i(_BoolToInt_2_i),
	.o(_BoolToInt_2_o)
);
BoolToInt BoolToInt_3(
	.clk(aclk),
	.i(_BoolToInt_3_i),
	.o(_BoolToInt_3_o)
);
BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_4 BitwiseIntConcat_3(
	.clk(aclk),
	.upper(_BitwiseIntConcat_3_upper),
	.lower(_BitwiseIntConcat_3_lower),
	.v(_BitwiseIntConcat_3_v)
);
always_ff @(posedge aclk) begin // state arvalid
	if(arvalid) if(arready) arvalid <= 1'b0;
	if(!arvalid) if(may_next_arvalid) arvalid <= 1'b1;
	if(_146) arvalid <= 1'b0;
end
always_ff @(posedge aclk) begin // state araddr
	if(!arvalid) if(may_next_arvalid) araddr <= _next_araddr_D0;
end
always_ff @(posedge aclk) begin // state arlen
	if(!arvalid) if(may_next_arvalid) arlen <= next_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = 3'd6;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _1;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _2;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _3;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = 1'd0;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = 1'd0;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rresp = 2'bxx;
	_rresp = rresp;
end
always_comb begin // combinatorial _rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rlast = 1'bx;
	_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_rlast = _rlast;
end
always_comb begin // combinatorial element_packet_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_packet_valid = 1'bx;
	element_packet_valid = 1'b0;
	if(rvalid) element_packet_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	element_packet_valid = element_packet_valid;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 16; _v0 = _v0 + 1) begin
if(rvalid) elements[_v0] = elements_2[_v0];
end
end
always_comb begin // combinatorial chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_offset = 4'dx;
	if(rvalid) chunk_offset = cur_chunk_align;
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 5'dx;
	if(rvalid) chunk_length = num_chunk_elements;
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(rvalid) last = is_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state num_in_flight
	num_in_flight <= _IntNarrow_4_out;
	if(_146) num_in_flight <= 1'd0;
end
always_ff @(posedge aclk) begin // state last_burst_in_flight
	if(!arvalid) if(may_next_arvalid) last_burst_in_flight <= _next_last_burst_in_flight_D0;
end
always_comb begin // combinatorial next_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_araddr = 64'dx;
	next_araddr = _BitwiseIntConcat_v;
end
always_comb begin // combinatorial _BitwiseIntConcat_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_upper = 58'dx;
	_BitwiseIntConcat_upper = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial _BitwiseIntConcat_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_lower = 6'dx;
	_BitwiseIntConcat_lower = 1'd0;
end
always_comb begin // combinatorial next_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_arlen = 6'dx;
	if(_chunks_are_left_D0) if(__23_D0) next_arlen = __26_D0;
	if(_chunks_are_left_D0) if(!__23_D0) next_arlen = _max_chunks_in_this_burst_D0;
end
always_comb begin // combinatorial next_last_burst_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_last_burst_in_flight = 1'bx;
	next_last_burst_in_flight = 1'b0;
	if(chunks_are_left) if(_23) next_last_burst_in_flight = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	next_last_burst_in_flight = next_last_burst_in_flight;
end
always_comb begin // combinatorial cur_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_burst_addr = 52'dx;
	cur_burst_addr = _BitwiseIntSplit_upper;
end
always_comb begin // combinatorial cur_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_align = 6'dx;
	cur_align = _BitwiseIntSplit_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_v = 58'dx;
	_BitwiseIntSplit_v = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial chunks_are_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunks_are_left = 1'bx;
	chunks_are_left = __14_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunks_are_left = chunks_are_left;
end
always_comb begin // combinatorial max_chunks_in_this_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	max_chunks_in_this_burst = 6'dx;
	if(chunks_are_left) max_chunks_in_this_burst = _18;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 17'dx;
	if(chunks_are_left) if(_23) _IntNarrow_in = __num_chunks_left_old_N1;
end
always_comb begin // combinatorial may_next_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_next_arvalid = 1'bx;
	may_next_arvalid = _39;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_next_arvalid = may_next_arvalid;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial next_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_burst_addr = 53'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) next_burst_addr = __45_D1;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_upper = 53'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_upper = next_burst_addr;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_lower = 6'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_lower = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_2_in = 59'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _IntNarrow_2_in = _BitwiseIntConcat_2_v;
end
always_comb begin // combinatorial _cur_start_chunk_addr_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_update = 1'bx;
	_cur_start_chunk_addr_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _cur_start_chunk_addr_update = 1'b1;
	if(request_new_burst) _cur_start_chunk_addr_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_update = _cur_start_chunk_addr_update;
end
always_comb begin // combinatorial _cur_start_chunk_addr_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_new = 58'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _cur_start_chunk_addr_new = _IntNarrow_2_out;
	if(_request_new_burst_D1) _cur_start_chunk_addr_new = _chunk_addr_D1;
end
always_comb begin // combinatorial next_num_chunks_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_num_chunks_left = 17'dx;
	if(!arvalid) if(may_next_arvalid) next_num_chunks_left = _IntNarrow_3_out;
end
always_comb begin // combinatorial _IntNarrow_3_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_3_in = 18'sdx;
	if(!arvalid) if(may_next_arvalid) _IntNarrow_3_in = _54;
end
always_comb begin // combinatorial _num_chunks_left_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_update = 1'bx;
	_num_chunks_left_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_update = 1'b1;
	if(request_new_burst) _num_chunks_left_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_update = _num_chunks_left_update;
end
always_comb begin // combinatorial _num_chunks_left_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_new = 17'dx;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_new = next_num_chunks_left;
	if(request_new_burst) _num_chunks_left_new = num_chunks;
end
always_comb begin // combinatorial _BoolToInt_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_i = 1'bx;
	_BoolToInt_i = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_i = _BoolToInt_i;
end
always_comb begin // combinatorial _Ternary_cond
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_cond = 1'bx;
	_Ternary_cond = _68;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Ternary_cond = _Ternary_cond;
end
always_comb begin // combinatorial _Ternary_a
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_a = 7'dx;
	_Ternary_a = _71;
end
always_comb begin // combinatorial _Ternary_b
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_b = 7'dx;
	_Ternary_b = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_4_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_4_in = 13'sdx;
	_IntNarrow_4_in = _73;
end
always_ff @(posedge aclk) begin // state final_chunk_align
	if(request_new_burst) final_chunk_align <= _BitwiseIntConcat_3_v;
end
always_ff @(posedge aclk) begin // state cur_chunk_align
	if(rvalid) cur_chunk_align <= 1'd0;
	if(request_new_burst) cur_chunk_align <= element_in_chunk_align;
end
always_comb begin // combinatorial elements_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_2 = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	if(rvalid) elements_2[0] = _75;
	if(rvalid) elements_2[1] = _76;
	if(rvalid) elements_2[2] = _77;
	if(rvalid) elements_2[3] = _78;
	if(rvalid) elements_2[4] = _79;
	if(rvalid) elements_2[5] = _80;
	if(rvalid) elements_2[6] = _81;
	if(rvalid) elements_2[7] = _82;
	if(rvalid) elements_2[8] = _83;
	if(rvalid) elements_2[9] = _84;
	if(rvalid) elements_2[10] = _85;
	if(rvalid) elements_2[11] = _86;
	if(rvalid) elements_2[12] = _87;
	if(rvalid) elements_2[13] = _88;
	if(rvalid) elements_2[14] = _89;
	if(rvalid) elements_2[15] = _90;
end
always_comb begin // combinatorial num_chunk_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunk_elements = 5'dx;
	if(rvalid) if(is_last) num_chunk_elements = _IntNarrow_5_out;
	if(rvalid) if(!is_last) num_chunk_elements = _101;
end
always_comb begin // combinatorial is_last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_last = 1'bx;
	if(rvalid) is_last = _95;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_last = is_last;
end
always_comb begin // combinatorial _IntNarrow_5_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_5_in = 6'sdx;
	if(rvalid) if(is_last) _IntNarrow_5_in = _99;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _113;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial chunk_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_addr = 58'dx;
	if(request_new_burst) chunk_addr = _BitwiseIntSplit_2_upper;
end
always_comb begin // combinatorial element_in_chunk_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_in_chunk_align = 4'dx;
	if(request_new_burst) element_in_chunk_align = _BitwiseIntSplit_2_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_2_v = 62'dx;
	if(request_new_burst) _BitwiseIntSplit_2_v = _115;
end
always_comb begin // combinatorial chunk_count_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_count_bits = 17'dx;
	if(request_new_burst) chunk_count_bits = _BitwiseIntSplit_3_upper;
end
always_comb begin // combinatorial final_alignment
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	final_alignment = 4'dx;
	if(request_new_burst) final_alignment = _BitwiseIntSplit_3_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_3_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_3_v = 21'dx;
	if(request_new_burst) _BitwiseIntSplit_3_v = _118;
end
always_comb begin // combinatorial num_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunks = 17'dx;
	if(request_new_burst) if(is_no_chunks) num_chunks = 1'd1;
	if(request_new_burst) if(!is_no_chunks) num_chunks = _128;
end
always_comb begin // combinatorial is_no_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_no_chunks = 1'bx;
	if(request_new_burst) is_no_chunks = _121;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_no_chunks = is_no_chunks;
end
always_comb begin // combinatorial _BoolToInt_2_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_2_i = 1'bx;
	if(request_new_burst) if(!is_no_chunks) _BoolToInt_2_i = _127;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_2_i = _BoolToInt_2_i;
end
always_comb begin // combinatorial _BoolToInt_3_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_3_i = 1'bx;
	if(request_new_burst) _BoolToInt_3_i = _138;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_3_i = _BoolToInt_3_i;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_upper = 1'dx;
	if(request_new_burst) _BitwiseIntConcat_3_upper = _BoolToInt_3_o;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BitwiseIntConcat_3_upper = _BitwiseIntConcat_3_upper;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_lower = 4'dx;
	if(request_new_burst) _BitwiseIntConcat_3_lower = final_alignment;
end
always_comb begin // combinatorial _cur_start_chunk_addr_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_rst = 1'bx;
	_cur_start_chunk_addr_rst = _142;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_rst = _cur_start_chunk_addr_rst;
end
always_comb begin // combinatorial _num_chunks_left_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_rst = 1'bx;
	_num_chunks_left_rst = _144;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_rst = _num_chunks_left_rst;
end
endmodule

// BitwiseIntConcat #(UPPER_TO: 2, LOWER_BITS: 4)
module BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_4(
	input clk,
	input wire[0:0] upper,
	input wire[3:0] lower,
	output /*mux_wire*/ logic[4:0] v
);

/*mux_wire*/ logic[4:0] v_bits;
/*mux_wire*/ logic[3:0] _UIntToBits_value;
wire[3:0] _UIntToBits_bits;
/*mux_wire*/ logic[0:0] _UIntToBits_2_value;
wire[0:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[4:0] _FromBits_bits;
wire[4:0] _FromBits_value;
UIntToBits_NUM_BITS_4 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_1 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_32 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 5'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 5'bxxxxx;
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
v_bits[4 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 4'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 1'dx;
	_UIntToBits_2_value = upper;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_UIntToBits_2_value = _UIntToBits_2_value;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 5'bxxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 32))
module FromBits_T_type_int_FROM_0_TO_32(
	input clk,
	input wire[4:0] bits,
	output /*mux_wire*/ logic[4:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 4)
module UIntToBits_NUM_BITS_4(
	input clk,
	input wire[3:0] value,
	output /*mux_wire*/ logic[3:0] bits
);

	assign bits = value;
endmodule

// BitwiseIntSplit #(TO: 1114127, LOWER_BITS: 4)
module BitwiseIntSplit_TO_1114127_LOWER_BITS_4(
	input clk,
	input wire[20:0] v,
	output /*mux_wire*/ logic[16:0] upper,
	output /*mux_wire*/ logic[3:0] lower
);

genvar _g0;
/*mux_wire*/ logic[20:0] v_bits;
/*mux_wire*/ logic[20:0] _UIntToBits_value;
wire[20:0] _UIntToBits_bits;
wire[3:0] _2;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_bits;
wire[3:0] _BitsToUInt_value;
wire[16:0] _3;
generate
for(_g0 = 0; _g0 < 17; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[4 + _g0];
end
endgenerate
/*mux_wire*/ logic[16:0] _FromBits_bits;
wire[16:0] _FromBits_value;
UIntToBits_NUM_BITS_21 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_4 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_69633 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 17'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 4'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 21'bxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 21'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 4'bxxxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 17'bxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 69633))
module FromBits_T_type_int_FROM_0_TO_69633(
	input clk,
	input wire[16:0] bits,
	output /*mux_wire*/ logic[16:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 21)
module UIntToBits_NUM_BITS_21(
	input clk,
	input wire[20:0] value,
	output /*mux_wire*/ logic[20:0] bits
);

	assign bits = value;
endmodule

// BitwiseIntSplit #(TO: 4611686018427387904, LOWER_BITS: 4)
module BitwiseIntSplit_TO_4611686018427387904_LOWER_BITS_4(
	input clk,
	input wire[61:0] v,
	output /*mux_wire*/ logic[57:0] upper,
	output /*mux_wire*/ logic[3:0] lower
);

genvar _g0;
/*mux_wire*/ logic[61:0] v_bits;
/*mux_wire*/ logic[61:0] _UIntToBits_value;
wire[61:0] _UIntToBits_bits;
wire[3:0] _2;
generate
for(_g0 = 0; _g0 < 4; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[3:0] _BitsToUInt_bits;
wire[3:0] _BitsToUInt_value;
wire[57:0] _3;
generate
for(_g0 = 0; _g0 < 58; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[4 + _g0];
end
endgenerate
/*mux_wire*/ logic[57:0] _FromBits_bits;
wire[57:0] _FromBits_value;
UIntToBits_NUM_BITS_62 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_4 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_288230376151711744 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 58'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 4'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 62'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 62'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 4'bxxxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 58'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 288230376151711744))
module FromBits_T_type_int_FROM_0_TO_288230376151711744(
	input clk,
	input wire[57:0] bits,
	output /*mux_wire*/ logic[57:0] value
);

assign value = bits;
endmodule

// BitsToUInt #(NUM_BITS: 4)
module BitsToUInt_NUM_BITS_4(
	input clk,
	input wire[3:0] bits,
	output /*mux_wire*/ logic[3:0] value
);

	assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 62)
module UIntToBits_NUM_BITS_62(
	input clk,
	input wire[61:0] value,
	output /*mux_wire*/ logic[61:0] bits
);

	assign bits = value;
endmodule

// IntNarrow #(FROM_I: -15, TO_I: 32, FROM: 0, TO: 17)
module IntNarrow_FROM_I_15_TO_I_32_FROM_0_TO_17(
	input clk,
	input wire signed[5:0] in,
	output /*mux_wire*/ logic[4:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: -1, TO_I: 3256, FROM: 0, TO: 3192)
module IntNarrow_FROM_I_1_TO_I_3256_FROM_0_TO_3192(
	input clk,
	input wire signed[12:0] in,
	output /*mux_wire*/ logic[11:0] out
);

	assign out = in;
endmodule

// Ternary #(T: type int #(FROM: 0, TO: 65))
module Ternary_T_type_int_FROM_0_TO_65(
	input clk,
	input wire cond,
	input wire[6:0] a,
	input wire[6:0] b,
	output /*mux_wire*/ logic[6:0] o
);

always_comb begin // combinatorial o
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	o = 7'dx;
	if(cond) o = a;
	if(!cond) o = b;
end
endmodule

// IntNarrow #(FROM_I: -64, TO_I: 69634, FROM: 0, TO: 69635)
module IntNarrow_FROM_I_64_TO_I_69634_FROM_0_TO_69635(
	input clk,
	input wire signed[17:0] in,
	output /*mux_wire*/ logic[16:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 288230376151711808, FROM: 0, TO: 288230376151711744)
module IntNarrow_FROM_I_0_TO_I_288230376151711808_FROM_0_TO_288230376151711744(
	input clk,
	input wire[58:0] in,
	output /*mux_wire*/ logic[57:0] out
);

	assign out = in;
endmodule

// BitwiseIntConcat #(UPPER_TO: 4503599627370497, LOWER_BITS: 6)
module BitwiseIntConcat_UPPER_TO_4503599627370497_LOWER_BITS_6(
	input clk,
	input wire[52:0] upper,
	input wire[5:0] lower,
	output /*mux_wire*/ logic[58:0] v
);

/*mux_wire*/ logic[58:0] v_bits;
/*mux_wire*/ logic[5:0] _UIntToBits_value;
wire[5:0] _UIntToBits_bits;
/*mux_wire*/ logic[52:0] _UIntToBits_2_value;
wire[52:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[58:0] _FromBits_bits;
wire[58:0] _FromBits_value;
UIntToBits_NUM_BITS_6 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_53 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_288230376151711808 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 59'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 59'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 53; _v0 = _v0 + 1) begin
v_bits[6 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 6'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 53'dx;
	_UIntToBits_2_value = upper;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 59'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 288230376151711808))
module FromBits_T_type_int_FROM_0_TO_288230376151711808(
	input clk,
	input wire[58:0] bits,
	output /*mux_wire*/ logic[58:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 53)
module UIntToBits_NUM_BITS_53(
	input clk,
	input wire[52:0] value,
	output /*mux_wire*/ logic[52:0] bits
);

	assign bits = value;
endmodule

// LatencyOffset #(T: type bool #(), OFFSET: 192)
module LatencyOffset_T_type_bool_OFFSET_192(
	input clk,
	input wire in,
	output /*mux_wire*/ logic out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 69635, FROM: 1, TO: 65)
module IntNarrow_FROM_I_0_TO_I_69635_FROM_1_TO_65(
	input clk,
	input wire[16:0] in,
	output /*mux_wire*/ logic[6:0] out
);

	assign out = in;
endmodule

// BitwiseIntSplit #(TO: 288230376151711744, LOWER_BITS: 6)
module BitwiseIntSplit_TO_288230376151711744_LOWER_BITS_6(
	input clk,
	input wire[57:0] v,
	output /*mux_wire*/ logic[51:0] upper,
	output /*mux_wire*/ logic[5:0] lower
);

genvar _g0;
/*mux_wire*/ logic[57:0] v_bits;
/*mux_wire*/ logic[57:0] _UIntToBits_value;
wire[57:0] _UIntToBits_bits;
wire[5:0] _2;
generate
for(_g0 = 0; _g0 < 6; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[5:0] _BitsToUInt_bits;
wire[5:0] _BitsToUInt_value;
wire[51:0] _3;
generate
for(_g0 = 0; _g0 < 52; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[6 + _g0];
end
endgenerate
/*mux_wire*/ logic[51:0] _FromBits_bits;
wire[51:0] _FromBits_value;
UIntToBits_NUM_BITS_58 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_6 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_4503599627370496 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 52'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 6'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 58'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 58'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 6'bxxxxxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 52'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 4503599627370496))
module FromBits_T_type_int_FROM_0_TO_4503599627370496(
	input clk,
	input wire[51:0] bits,
	output /*mux_wire*/ logic[51:0] value
);

assign value = bits;
endmodule

// BitsToUInt #(NUM_BITS: 6)
module BitsToUInt_NUM_BITS_6(
	input clk,
	input wire[5:0] bits,
	output /*mux_wire*/ logic[5:0] value
);

	assign value = bits;
endmodule

// BitwiseIntConcat #(UPPER_TO: 288230376151711744, LOWER_BITS: 6)
module BitwiseIntConcat_UPPER_TO_288230376151711744_LOWER_BITS_6(
	input clk,
	input wire[57:0] upper,
	input wire[5:0] lower,
	output /*mux_wire*/ logic[63:0] v
);

/*mux_wire*/ logic[63:0] v_bits;
/*mux_wire*/ logic[5:0] _UIntToBits_value;
wire[5:0] _UIntToBits_bits;
/*mux_wire*/ logic[57:0] _UIntToBits_2_value;
wire[57:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[63:0] _FromBits_bits;
wire[63:0] _FromBits_value;
UIntToBits_NUM_BITS_6 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_58 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_18446744073709551616 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 64'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 6; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 58; _v0 = _v0 + 1) begin
v_bits[6 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 6'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 58'dx;
	_UIntToBits_2_value = upper;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// UIntToBits #(NUM_BITS: 58)
module UIntToBits_NUM_BITS_58(
	input clk,
	input wire[57:0] value,
	output /*mux_wire*/ logic[57:0] bits
);

	assign bits = value;
endmodule

// UIntToBits #(NUM_BITS: 6)
module UIntToBits_NUM_BITS_6(
	input clk,
	input wire[5:0] value,
	output /*mux_wire*/ logic[5:0] bits
);

	assign bits = value;
endmodule

// SlowState #(T: type int #(FROM: 0, TO: 69635), RESET_TO: 0, OLD_DELAY: 2, NEW_DELAY: 0)
module SlowState_T_type_int_FROM_0_TO_69635_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0(
	input clk,
	input wire rst,
	output /*state*/ logic[16:0] old,
	output /*mux_wire*/ logic may_update,
	input wire update,
	input wire[16:0] new_1
);

genvar _g0;
/*mux_wire*/ logic _cross_rst_in;
/*mux_wire*/ logic[16:0] new_s;
/*mux_wire*/ logic update_s;
/*mux_wire*/ logic update_old;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
/*mux_wire*/ logic[16:0] new_old;
/*mux_wire*/ logic[16:0] _LatencyOffset_2_in;
wire[16:0] _LatencyOffset_2_out;
wire _cross_rst_out;
/*latency*/ logic __cross_rst_out_N1; always_ff @(posedge clk) begin __cross_rst_out_N1 <= _cross_rst_out; end
/*latency*/ logic __cross_rst_out_D0; always_ff @(posedge clk) begin __cross_rst_out_D0 <= __cross_rst_out_N1; end
/*state*/ logic[1:0] cooldown;
wire _8 = cooldown[0];
wire _11;
assign _11 = update_s | __cross_rst_out_D0;
/*mux_wire*/ logic _Repeat_v;
wire[1:0] _Repeat_result;
wire[0:0] _12;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _12[_g0] = cooldown[1 + _g0];
end
endgenerate
CrossDomain_T_type_bool cross_rst(
	.in_clk(clk),
	.in(_cross_rst_in),
	.out(_cross_rst_out)
);
LatencyOffset_T_type_bool_OFFSET_2 LatencyOffset(
	.clk(clk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
LatencyOffset_T_type_int_FROM_0_TO_69635_OFFSET_2 LatencyOffset_2(
	.clk(clk),
	.in(_LatencyOffset_2_in),
	.out(_LatencyOffset_2_out)
);
Repeat_T_type_bool_SIZE_2 Repeat(
	.clk(clk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
always_comb begin // combinatorial _cross_rst_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_rst_in = 1'bx;
	_cross_rst_in = rst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_rst_in = _cross_rst_in;
end
always_ff @(posedge clk) begin // state old
	if(_cross_rst_out) old <= 17'd0;
	if(!_cross_rst_out) if(update_old) old <= new_old;
end
always_comb begin // combinatorial new_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_s = 17'dx;
	if(update) new_s = new_1;
end
always_comb begin // combinatorial update_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_s = 1'bx;
	if(update) update_s = 1'b1;
	if(!update) update_s = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_s = update_s;
end
always_comb begin // combinatorial update_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_old = 1'bx;
	update_old = _LatencyOffset_out;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_old = update_old;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = update_s;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial new_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_old = 17'dx;
	new_old = _LatencyOffset_2_out;
end
always_comb begin // combinatorial _LatencyOffset_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_2_in = 17'dx;
	_LatencyOffset_2_in = new_s;
end
always_comb begin // combinatorial may_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_update = 1'bx;
	may_update = _8;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_update = may_update;
end
always_ff @(posedge clk) begin // state cooldown
	if(_11) cooldown <= _Repeat_result;
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(!_11) cooldown[_v0] <= _12[_v0];
end
	if(!_11) cooldown[1] <= 1'b1;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	if(_11) _Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
endmodule

// LatencyOffset #(T: type int #(FROM: 0, TO: 69635), OFFSET: -2)
module LatencyOffset_T_type_int_FROM_0_TO_69635_OFFSET_2(
	input clk,
	input wire[16:0] in,
	output /*mux_wire*/ logic[16:0] out
);

	assign out = in;
endmodule

// SlowState #(T: type int #(FROM: 0, TO: 288230376151711744), RESET_TO: 0, OLD_DELAY: 1, NEW_DELAY: 1)
module SlowState_T_type_int_FROM_0_TO_288230376151711744_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1(
	input clk,
	input wire rst,
	output /*state*/ logic[57:0] old,
	output /*mux_wire*/ logic may_update,
	input wire update,
	input wire[57:0] new_1
);

/*latency*/ logic _update_D1; always_ff @(posedge clk) begin _update_D1 <= update; end
genvar _g0;
/*mux_wire*/ logic _cross_rst_in;
/*mux_wire*/ logic[57:0] new_s;
/*mux_wire*/ logic update_s;
/*mux_wire*/ logic update_old;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
/*latency*/ logic __LatencyOffset_out_N1; always_ff @(posedge clk) begin __LatencyOffset_out_N1 <= _LatencyOffset_out; end
/*mux_wire*/ logic[57:0] new_old;
/*mux_wire*/ logic[57:0] _LatencyOffset_2_in;
wire[57:0] _LatencyOffset_2_out;
wire _cross_rst_out;
/*latency*/ logic __cross_rst_out_D0; always_ff @(posedge clk) begin __cross_rst_out_D0 <= _cross_rst_out; end
/*state*/ logic[1:0] cooldown;
wire _8 = cooldown[0];
wire _11;
assign _11 = update_s | __cross_rst_out_D0;
/*mux_wire*/ logic _Repeat_v;
wire[1:0] _Repeat_result;
wire[0:0] _12;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _12[_g0] = cooldown[1 + _g0];
end
endgenerate
CrossDomain_T_type_bool cross_rst(
	.in_clk(clk),
	.in(_cross_rst_in),
	.out(_cross_rst_out)
);
LatencyOffset_T_type_bool_OFFSET_2 LatencyOffset(
	.clk(clk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
LatencyOffset_T_type_int_FROM_0_TO_288230376151711744_OFFSET_2 LatencyOffset_2(
	.clk(clk),
	.in(_LatencyOffset_2_in),
	.out(_LatencyOffset_2_out)
);
Repeat_T_type_bool_SIZE_2 Repeat(
	.clk(clk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
always_comb begin // combinatorial _cross_rst_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_rst_in = 1'bx;
	_cross_rst_in = rst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_rst_in = _cross_rst_in;
end
always_ff @(posedge clk) begin // state old
	if(_cross_rst_out) old <= 58'd0;
	if(!_cross_rst_out) if(update_old) old <= new_old;
end
always_comb begin // combinatorial new_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_s = 58'dx;
	if(_update_D1) new_s = new_1;
end
always_comb begin // combinatorial update_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_s = 1'bx;
	if(update) update_s = 1'b1;
	if(!update) update_s = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_s = update_s;
end
always_comb begin // combinatorial update_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_old = 1'bx;
	update_old = __LatencyOffset_out_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_old = update_old;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = update_s;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial new_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_old = 58'dx;
	new_old = _LatencyOffset_2_out;
end
always_comb begin // combinatorial _LatencyOffset_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_2_in = 58'dx;
	_LatencyOffset_2_in = new_s;
end
always_comb begin // combinatorial may_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_update = 1'bx;
	may_update = _8;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_update = may_update;
end
always_ff @(posedge clk) begin // state cooldown
	if(_11) cooldown <= _Repeat_result;
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(!_11) cooldown[_v0] <= _12[_v0];
end
	if(!_11) cooldown[1] <= 1'b1;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	if(_11) _Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
endmodule

// LatencyOffset #(T: type int #(FROM: 0, TO: 288230376151711744), OFFSET: -2)
module LatencyOffset_T_type_int_FROM_0_TO_288230376151711744_OFFSET_2(
	input clk,
	input wire[57:0] in,
	output /*mux_wire*/ logic[57:0] out
);

	assign out = in;
endmodule

// axi_array_burst_reader #(AXI_WIDTH: 64, ADDR_ALIGN: 2, COUNT_TO: 65536, ATO: 18446744073709551616)
module axi_array_burst_reader_AXI_WIDTH_64_ADDR_ALIGN_2_COUNT_TO_65536_ATO_18446744073709551616(
	input aclk,
	input wire aresetn,
	output /*state*/ logic arvalid,
	input wire arready,
	output /*state*/ logic[63:0] araddr,
	output /*state*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[63:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire is_ready_to_receive_lots_of_data,
	output /*mux_wire*/ logic element_packet_valid,
	output /*mux_wire*/ logic[15:0] elements[3:0],
	output /*mux_wire*/ logic[1:0] chunk_offset,
	output /*mux_wire*/ logic[2:0] chunk_length,
	output /*mux_wire*/ logic last,
	input wire[10:0] max_in_flight,
	output /*mux_wire*/ logic may_request_new_burst,
	input wire request_new_burst,
	input wire[63:0] start_addr,
	input wire[15:0] count
);

/*latency*/ logic _arvalid_D1; always_ff @(posedge aclk) begin _arvalid_D1 <= arvalid; end
/*latency*/ logic _request_new_burst_D1; always_ff @(posedge aclk) begin _request_new_burst_D1 <= request_new_burst; end
genvar _g0;
localparam[1:0] _1 = 2'b01;
localparam[2:0] _2 = 3'b000;
localparam[3:0] _3 = 4'b0010;
/*mux_wire*/ logic[1:0] _rresp;
/*mux_wire*/ logic _rlast;
/*state*/ logic[11:0] num_in_flight;
/*state*/ logic last_burst_in_flight;
/*mux_wire*/ logic[63:0] next_araddr;
/*latency*/ logic[63:0] _next_araddr_D0; always_ff @(posedge aclk) begin _next_araddr_D0 <= next_araddr; end
wire[60:0] _cur_start_chunk_addr_old;
/*mux_wire*/ logic[60:0] _BitwiseIntConcat_upper;
/*mux_wire*/ logic[2:0] _BitwiseIntConcat_lower;
wire[63:0] _BitwiseIntConcat_v;
/*mux_wire*/ logic[7:0] next_arlen;
/*mux_wire*/ logic next_last_burst_in_flight;
/*latency*/ logic _next_last_burst_in_flight_D0; always_ff @(posedge aclk) begin _next_last_burst_in_flight_D0 <= next_last_burst_in_flight; end
/*mux_wire*/ logic[52:0] cur_burst_addr;
/*mux_wire*/ logic[7:0] cur_align;
/*mux_wire*/ logic[60:0] _BitwiseIntSplit_v;
wire[52:0] _BitwiseIntSplit_upper;
wire[7:0] _BitwiseIntSplit_lower;
/*mux_wire*/ logic chunks_are_left;
/*latency*/ logic _chunks_are_left_D0; always_ff @(posedge aclk) begin _chunks_are_left_D0 <= chunks_are_left; end
wire[14:0] _num_chunks_left_old;
/*latency*/ logic[14:0] __num_chunks_left_old_N1; always_ff @(posedge aclk) begin __num_chunks_left_old_N1 <= _num_chunks_left_old; end
/*latency*/ logic[14:0] __num_chunks_left_old_D0; always_ff @(posedge aclk) begin __num_chunks_left_old_D0 <= __num_chunks_left_old_N1; end
wire _14;
assign _14 = _num_chunks_left_old > 1'd0;
/*latency*/ logic __14_N1; always_ff @(posedge aclk) begin __14_N1 <= _14; end
/*mux_wire*/ logic[7:0] max_chunks_in_this_burst;
/*latency*/ logic[7:0] _max_chunks_in_this_burst_D0; always_ff @(posedge aclk) begin _max_chunks_in_this_burst_D0 <= max_chunks_in_this_burst; end
wire[7:0] _18;
assign _18 = 8'd255 - cur_align;
wire[8:0] _22;
assign _22 = max_chunks_in_this_burst + 1'd1;
wire _23;
assign _23 = __num_chunks_left_old_N1 <= _22;
/*latency*/ logic __23_D0; always_ff @(posedge aclk) begin __23_D0 <= _23; end
/*mux_wire*/ logic[14:0] _IntNarrow_in;
wire[8:0] _IntNarrow_out;
wire[7:0] _26;
assign _26 = _IntNarrow_out - 1'd1;
/*latency*/ logic[7:0] __26_D0; always_ff @(posedge aclk) begin __26_D0 <= _26; end
/*mux_wire*/ logic may_next_arvalid;
/*latency*/ logic _may_next_arvalid_D1; always_ff @(posedge aclk) begin _may_next_arvalid_D1 <= may_next_arvalid; end
wire _num_chunks_left_may_update;
wire _30;
assign _30 = _chunks_are_left_D0 & _num_chunks_left_may_update;
wire _cur_start_chunk_addr_may_update;
wire _32;
assign _32 = _30 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
wire _34;
assign _34 = _32 & _LatencyOffset_out;
wire signed[11:0] _37;
assign _37 = max_in_flight - 9'd256;
wire _38;
assign _38 = $signed({1'b0, num_in_flight}) <= _37;
wire _39;
assign _39 = _34 & _38;
/*mux_wire*/ logic[53:0] next_burst_addr;
wire[53:0] _45;
assign _45 = cur_burst_addr + 1'd1;
/*latency*/ logic[53:0] __45_D0; always_ff @(posedge aclk) begin __45_D0 <= _45; end
/*latency*/ logic[53:0] __45_D1; always_ff @(posedge aclk) begin __45_D1 <= __45_D0; end
/*mux_wire*/ logic[53:0] _BitwiseIntConcat_2_upper;
/*mux_wire*/ logic[7:0] _BitwiseIntConcat_2_lower;
wire[61:0] _BitwiseIntConcat_2_v;
/*mux_wire*/ logic[61:0] _IntNarrow_2_in;
wire[60:0] _IntNarrow_2_out;
/*mux_wire*/ logic _cur_start_chunk_addr_update;
/*mux_wire*/ logic[60:0] _cur_start_chunk_addr_new;
/*mux_wire*/ logic[14:0] next_num_chunks_left;
wire[8:0] _53;
assign _53 = next_arlen + 1'd1;
wire signed[15:0] _54;
assign _54 = __num_chunks_left_old_D0 - _53;
/*mux_wire*/ logic signed[15:0] _IntNarrow_3_in;
wire[14:0] _IntNarrow_3_out;
/*mux_wire*/ logic _num_chunks_left_update;
/*mux_wire*/ logic[14:0] _num_chunks_left_new;
/*mux_wire*/ logic _BoolToInt_i;
wire[0:0] _BoolToInt_o;
wire signed[12:0] _64;
assign _64 = num_in_flight - _BoolToInt_o;
wire _66;
assign _66 = !arvalid;
wire _68;
assign _68 = _66 & may_next_arvalid;
wire[8:0] _71;
assign _71 = next_arlen + 1'd1;
/*mux_wire*/ logic _Ternary_cond;
/*mux_wire*/ logic[8:0] _Ternary_a;
/*mux_wire*/ logic[8:0] _Ternary_b;
wire[8:0] _Ternary_o;
wire signed[12:0] _73;
assign _73 = _64 + $signed({1'b0, _Ternary_o});
/*mux_wire*/ logic signed[12:0] _IntNarrow_4_in;
wire[11:0] _IntNarrow_4_out;
/*state*/ logic[2:0] final_chunk_align;
/*state*/ logic[1:0] cur_chunk_align;
/*mux_wire*/ logic[15:0] elements_2[3:0];
wire[15:0] _75;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _75[_g0] = rdata[_g0];
end
endgenerate
wire[15:0] _76;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _76[_g0] = rdata[16 + _g0];
end
endgenerate
wire[15:0] _77;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _77[_g0] = rdata[32 + _g0];
end
endgenerate
wire[15:0] _78;
generate
for(_g0 = 0; _g0 < 16; _g0 = _g0 + 1) begin
assign _78[_g0] = rdata[48 + _g0];
end
endgenerate
/*mux_wire*/ logic[2:0] num_chunk_elements;
/*mux_wire*/ logic is_last;
wire _81;
assign _81 = num_in_flight == 1'd1;
wire _83;
assign _83 = _81 & last_burst_in_flight;
wire signed[3:0] _87;
assign _87 = final_chunk_align - cur_chunk_align;
/*mux_wire*/ logic signed[3:0] _IntNarrow_5_in;
wire[2:0] _IntNarrow_5_out;
wire[2:0] _89;
assign _89 = 3'd4 - cur_chunk_align;
wire _97;
assign _97 = !chunks_are_left;
/*latency*/ logic __97_D0; always_ff @(posedge aclk) begin __97_D0 <= _97; end
wire _99;
assign _99 = __97_D0 & _num_chunks_left_may_update;
wire _101;
assign _101 = _99 & _cur_start_chunk_addr_may_update;
/*mux_wire*/ logic[60:0] chunk_addr;
/*latency*/ logic[60:0] _chunk_addr_D1; always_ff @(posedge aclk) begin _chunk_addr_D1 <= chunk_addr; end
/*mux_wire*/ logic[1:0] element_in_chunk_align;
wire[62:0] _103;
assign _103 = start_addr / 2'd2;
/*mux_wire*/ logic[62:0] _BitwiseIntSplit_2_v;
wire[60:0] _BitwiseIntSplit_2_upper;
wire[1:0] _BitwiseIntSplit_2_lower;
/*mux_wire*/ logic[14:0] chunk_count_bits;
/*mux_wire*/ logic[1:0] final_alignment;
wire[16:0] _106;
assign _106 = count + element_in_chunk_align;
/*mux_wire*/ logic[16:0] _BitwiseIntSplit_3_v;
wire[14:0] _BitwiseIntSplit_3_upper;
wire[1:0] _BitwiseIntSplit_3_lower;
/*mux_wire*/ logic[14:0] num_chunks;
/*mux_wire*/ logic is_no_chunks;
wire _109;
assign _109 = chunk_count_bits == 1'd0;
wire _115;
assign _115 = final_alignment != 1'd0;
/*mux_wire*/ logic _BoolToInt_2_i;
wire[0:0] _BoolToInt_2_o;
wire[14:0] _116;
assign _116 = chunk_count_bits + _BoolToInt_2_o;
wire _122;
assign _122 = !is_no_chunks;
wire _125;
assign _125 = final_alignment == 1'd0;
wire _126;
assign _126 = _122 & _125;
/*mux_wire*/ logic _BoolToInt_3_i;
wire[0:0] _BoolToInt_3_o;
/*mux_wire*/ logic[0:0] _BitwiseIntConcat_3_upper;
/*mux_wire*/ logic[1:0] _BitwiseIntConcat_3_lower;
wire[2:0] _BitwiseIntConcat_3_v;
wire _130;
assign _130 = !aresetn;
/*mux_wire*/ logic _cur_start_chunk_addr_rst;
wire _132;
assign _132 = !aresetn;
/*mux_wire*/ logic _num_chunks_left_rst;
wire _134;
assign _134 = !aresetn;
SlowState_T_type_int_FROM_0_TO_2305843009213693952_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1 cur_start_chunk_addr(
	.clk(aclk),
	.rst(_cur_start_chunk_addr_rst),
	.old(_cur_start_chunk_addr_old),
	.may_update(_cur_start_chunk_addr_may_update),
	.update(_cur_start_chunk_addr_update),
	.new_1(_cur_start_chunk_addr_new)
);
SlowState_T_type_int_FROM_0_TO_16387_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0 num_chunks_left(
	.clk(aclk),
	.rst(_num_chunks_left_rst),
	.old(_num_chunks_left_old),
	.may_update(_num_chunks_left_may_update),
	.update(_num_chunks_left_update),
	.new_1(_num_chunks_left_new)
);
BitwiseIntConcat_UPPER_TO_2305843009213693952_LOWER_BITS_3 BitwiseIntConcat(
	.clk(aclk),
	.upper(_BitwiseIntConcat_upper),
	.lower(_BitwiseIntConcat_lower),
	.v(_BitwiseIntConcat_v)
);
BitwiseIntSplit_TO_2305843009213693952_LOWER_BITS_8 BitwiseIntSplit(
	.clk(aclk),
	.v(_BitwiseIntSplit_v),
	.upper(_BitwiseIntSplit_upper),
	.lower(_BitwiseIntSplit_lower)
);
IntNarrow_FROM_I_0_TO_I_16387_FROM_1_TO_257 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
LatencyOffset_T_type_bool_OFFSET_384 LatencyOffset(
	.clk(aclk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
BitwiseIntConcat_UPPER_TO_9007199254740993_LOWER_BITS_8 BitwiseIntConcat_2(
	.clk(aclk),
	.upper(_BitwiseIntConcat_2_upper),
	.lower(_BitwiseIntConcat_2_lower),
	.v(_BitwiseIntConcat_2_v)
);
IntNarrow_FROM_I_0_TO_I_2305843009213694208_FROM_0_TO_2305843009213693952 IntNarrow_2(
	.clk(aclk),
	.in(_IntNarrow_2_in),
	.out(_IntNarrow_2_out)
);
IntNarrow_FROM_I_256_TO_I_16386_FROM_0_TO_16387 IntNarrow_3(
	.clk(aclk),
	.in(_IntNarrow_3_in),
	.out(_IntNarrow_3_out)
);
BoolToInt BoolToInt(
	.clk(aclk),
	.i(_BoolToInt_i),
	.o(_BoolToInt_o)
);
Ternary_T_type_int_FROM_0_TO_257 Ternary(
	.clk(aclk),
	.cond(_Ternary_cond),
	.a(_Ternary_a),
	.b(_Ternary_b),
	.o(_Ternary_o)
);
IntNarrow_FROM_I_1_TO_I_3640_FROM_0_TO_3384 IntNarrow_4(
	.clk(aclk),
	.in(_IntNarrow_4_in),
	.out(_IntNarrow_4_out)
);
IntNarrow_FROM_I_3_TO_I_8_FROM_0_TO_5 IntNarrow_5(
	.clk(aclk),
	.in(_IntNarrow_5_in),
	.out(_IntNarrow_5_out)
);
BitwiseIntSplit_TO_9223372036854775808_LOWER_BITS_2 BitwiseIntSplit_2(
	.clk(aclk),
	.v(_BitwiseIntSplit_2_v),
	.upper(_BitwiseIntSplit_2_upper),
	.lower(_BitwiseIntSplit_2_lower)
);
BitwiseIntSplit_TO_65539_LOWER_BITS_2 BitwiseIntSplit_3(
	.clk(aclk),
	.v(_BitwiseIntSplit_3_v),
	.upper(_BitwiseIntSplit_3_upper),
	.lower(_BitwiseIntSplit_3_lower)
);
BoolToInt BoolToInt_2(
	.clk(aclk),
	.i(_BoolToInt_2_i),
	.o(_BoolToInt_2_o)
);
BoolToInt BoolToInt_3(
	.clk(aclk),
	.i(_BoolToInt_3_i),
	.o(_BoolToInt_3_o)
);
BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_2 BitwiseIntConcat_3(
	.clk(aclk),
	.upper(_BitwiseIntConcat_3_upper),
	.lower(_BitwiseIntConcat_3_lower),
	.v(_BitwiseIntConcat_3_v)
);
always_ff @(posedge aclk) begin // state arvalid
	if(arvalid) if(arready) arvalid <= 1'b0;
	if(!arvalid) if(may_next_arvalid) arvalid <= 1'b1;
	if(_134) arvalid <= 1'b0;
end
always_ff @(posedge aclk) begin // state araddr
	if(!arvalid) if(may_next_arvalid) araddr <= _next_araddr_D0;
end
always_ff @(posedge aclk) begin // state arlen
	if(!arvalid) if(may_next_arvalid) arlen <= next_arlen;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = 2'd3;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _1;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _2;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _3;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = 1'd0;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = 1'd0;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rresp = 2'bxx;
	_rresp = rresp;
end
always_comb begin // combinatorial _rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rlast = 1'bx;
	_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_rlast = _rlast;
end
always_comb begin // combinatorial element_packet_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_packet_valid = 1'bx;
	element_packet_valid = 1'b0;
	if(rvalid) element_packet_valid = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	element_packet_valid = element_packet_valid;
end
always_comb begin // combinatorial elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements = '{16'bxxxxxxxxxxxxxxxx, 16'bxxxxxxxxxxxxxxxx, 16'bxxxxxxxxxxxxxxxx, 16'bxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 4; _v0 = _v0 + 1) begin
if(rvalid) elements[_v0] = elements_2[_v0];
end
end
always_comb begin // combinatorial chunk_offset
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_offset = 2'dx;
	if(rvalid) chunk_offset = cur_chunk_align;
end
always_comb begin // combinatorial chunk_length
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_length = 3'dx;
	if(rvalid) chunk_length = num_chunk_elements;
end
always_comb begin // combinatorial last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	last = 1'bx;
	if(rvalid) last = is_last;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	last = last;
end
always_ff @(posedge aclk) begin // state num_in_flight
	num_in_flight <= _IntNarrow_4_out;
	if(_134) num_in_flight <= 1'd0;
end
always_ff @(posedge aclk) begin // state last_burst_in_flight
	if(!arvalid) if(may_next_arvalid) last_burst_in_flight <= _next_last_burst_in_flight_D0;
end
always_comb begin // combinatorial next_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_araddr = 64'dx;
	next_araddr = _BitwiseIntConcat_v;
end
always_comb begin // combinatorial _BitwiseIntConcat_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_upper = 61'dx;
	_BitwiseIntConcat_upper = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial _BitwiseIntConcat_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_lower = 3'dx;
	_BitwiseIntConcat_lower = 1'd0;
end
always_comb begin // combinatorial next_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_arlen = 8'dx;
	if(_chunks_are_left_D0) if(__23_D0) next_arlen = __26_D0;
	if(_chunks_are_left_D0) if(!__23_D0) next_arlen = _max_chunks_in_this_burst_D0;
end
always_comb begin // combinatorial next_last_burst_in_flight
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_last_burst_in_flight = 1'bx;
	next_last_burst_in_flight = 1'b0;
	if(chunks_are_left) if(_23) next_last_burst_in_flight = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	next_last_burst_in_flight = next_last_burst_in_flight;
end
always_comb begin // combinatorial cur_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_burst_addr = 53'dx;
	cur_burst_addr = _BitwiseIntSplit_upper;
end
always_comb begin // combinatorial cur_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	cur_align = 8'dx;
	cur_align = _BitwiseIntSplit_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_v = 61'dx;
	_BitwiseIntSplit_v = _cur_start_chunk_addr_old;
end
always_comb begin // combinatorial chunks_are_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunks_are_left = 1'bx;
	chunks_are_left = __14_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	chunks_are_left = chunks_are_left;
end
always_comb begin // combinatorial max_chunks_in_this_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	max_chunks_in_this_burst = 8'dx;
	if(chunks_are_left) max_chunks_in_this_burst = _18;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 15'dx;
	if(chunks_are_left) if(_23) _IntNarrow_in = __num_chunks_left_old_N1;
end
always_comb begin // combinatorial may_next_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_next_arvalid = 1'bx;
	may_next_arvalid = _39;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_next_arvalid = may_next_arvalid;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = is_ready_to_receive_lots_of_data;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial next_burst_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_burst_addr = 54'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) next_burst_addr = __45_D1;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_upper = 54'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_upper = next_burst_addr;
end
always_comb begin // combinatorial _BitwiseIntConcat_2_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_2_lower = 8'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _BitwiseIntConcat_2_lower = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_2_in = 62'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _IntNarrow_2_in = _BitwiseIntConcat_2_v;
end
always_comb begin // combinatorial _cur_start_chunk_addr_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_update = 1'bx;
	_cur_start_chunk_addr_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _cur_start_chunk_addr_update = 1'b1;
	if(request_new_burst) _cur_start_chunk_addr_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_update = _cur_start_chunk_addr_update;
end
always_comb begin // combinatorial _cur_start_chunk_addr_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_new = 61'dx;
	if(!_arvalid_D1) if(_may_next_arvalid_D1) _cur_start_chunk_addr_new = _IntNarrow_2_out;
	if(_request_new_burst_D1) _cur_start_chunk_addr_new = _chunk_addr_D1;
end
always_comb begin // combinatorial next_num_chunks_left
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	next_num_chunks_left = 15'dx;
	if(!arvalid) if(may_next_arvalid) next_num_chunks_left = _IntNarrow_3_out;
end
always_comb begin // combinatorial _IntNarrow_3_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_3_in = 16'sdx;
	if(!arvalid) if(may_next_arvalid) _IntNarrow_3_in = _54;
end
always_comb begin // combinatorial _num_chunks_left_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_update = 1'bx;
	_num_chunks_left_update = 1'b0;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_update = 1'b1;
	if(request_new_burst) _num_chunks_left_update = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_update = _num_chunks_left_update;
end
always_comb begin // combinatorial _num_chunks_left_new
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_new = 15'dx;
	if(!arvalid) if(may_next_arvalid) _num_chunks_left_new = next_num_chunks_left;
	if(request_new_burst) _num_chunks_left_new = num_chunks;
end
always_comb begin // combinatorial _BoolToInt_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_i = 1'bx;
	_BoolToInt_i = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_i = _BoolToInt_i;
end
always_comb begin // combinatorial _Ternary_cond
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_cond = 1'bx;
	_Ternary_cond = _68;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Ternary_cond = _Ternary_cond;
end
always_comb begin // combinatorial _Ternary_a
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_a = 9'dx;
	_Ternary_a = _71;
end
always_comb begin // combinatorial _Ternary_b
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Ternary_b = 9'dx;
	_Ternary_b = 1'd0;
end
always_comb begin // combinatorial _IntNarrow_4_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_4_in = 13'sdx;
	_IntNarrow_4_in = _73;
end
always_ff @(posedge aclk) begin // state final_chunk_align
	if(request_new_burst) final_chunk_align <= _BitwiseIntConcat_3_v;
end
always_ff @(posedge aclk) begin // state cur_chunk_align
	if(rvalid) cur_chunk_align <= 1'd0;
	if(request_new_burst) cur_chunk_align <= element_in_chunk_align;
end
always_comb begin // combinatorial elements_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	elements_2 = '{16'bxxxxxxxxxxxxxxxx, 16'bxxxxxxxxxxxxxxxx, 16'bxxxxxxxxxxxxxxxx, 16'bxxxxxxxxxxxxxxxx};
	if(rvalid) elements_2[0] = _75;
	if(rvalid) elements_2[1] = _76;
	if(rvalid) elements_2[2] = _77;
	if(rvalid) elements_2[3] = _78;
end
always_comb begin // combinatorial num_chunk_elements
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunk_elements = 3'dx;
	if(rvalid) if(is_last) num_chunk_elements = _IntNarrow_5_out;
	if(rvalid) if(!is_last) num_chunk_elements = _89;
end
always_comb begin // combinatorial is_last
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_last = 1'bx;
	if(rvalid) is_last = _83;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_last = is_last;
end
always_comb begin // combinatorial _IntNarrow_5_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_5_in = 4'sdx;
	if(rvalid) if(is_last) _IntNarrow_5_in = _87;
end
always_comb begin // combinatorial may_request_new_burst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_request_new_burst = 1'bx;
	may_request_new_burst = _101;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_request_new_burst = may_request_new_burst;
end
always_comb begin // combinatorial chunk_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_addr = 61'dx;
	if(request_new_burst) chunk_addr = _BitwiseIntSplit_2_upper;
end
always_comb begin // combinatorial element_in_chunk_align
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	element_in_chunk_align = 2'dx;
	if(request_new_burst) element_in_chunk_align = _BitwiseIntSplit_2_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_2_v = 63'dx;
	if(request_new_burst) _BitwiseIntSplit_2_v = _103;
end
always_comb begin // combinatorial chunk_count_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	chunk_count_bits = 15'dx;
	if(request_new_burst) chunk_count_bits = _BitwiseIntSplit_3_upper;
end
always_comb begin // combinatorial final_alignment
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	final_alignment = 2'dx;
	if(request_new_burst) final_alignment = _BitwiseIntSplit_3_lower;
end
always_comb begin // combinatorial _BitwiseIntSplit_3_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntSplit_3_v = 17'dx;
	if(request_new_burst) _BitwiseIntSplit_3_v = _106;
end
always_comb begin // combinatorial num_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	num_chunks = 15'dx;
	if(request_new_burst) if(is_no_chunks) num_chunks = 1'd1;
	if(request_new_burst) if(!is_no_chunks) num_chunks = _116;
end
always_comb begin // combinatorial is_no_chunks
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	is_no_chunks = 1'bx;
	if(request_new_burst) is_no_chunks = _109;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	is_no_chunks = is_no_chunks;
end
always_comb begin // combinatorial _BoolToInt_2_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_2_i = 1'bx;
	if(request_new_burst) if(!is_no_chunks) _BoolToInt_2_i = _115;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_2_i = _BoolToInt_2_i;
end
always_comb begin // combinatorial _BoolToInt_3_i
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BoolToInt_3_i = 1'bx;
	if(request_new_burst) _BoolToInt_3_i = _126;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BoolToInt_3_i = _BoolToInt_3_i;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_upper = 1'dx;
	if(request_new_burst) _BitwiseIntConcat_3_upper = _BoolToInt_3_o;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_BitwiseIntConcat_3_upper = _BitwiseIntConcat_3_upper;
end
always_comb begin // combinatorial _BitwiseIntConcat_3_lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitwiseIntConcat_3_lower = 2'dx;
	if(request_new_burst) _BitwiseIntConcat_3_lower = final_alignment;
end
always_comb begin // combinatorial _cur_start_chunk_addr_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cur_start_chunk_addr_rst = 1'bx;
	_cur_start_chunk_addr_rst = _130;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cur_start_chunk_addr_rst = _cur_start_chunk_addr_rst;
end
always_comb begin // combinatorial _num_chunks_left_rst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_num_chunks_left_rst = 1'bx;
	_num_chunks_left_rst = _132;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_num_chunks_left_rst = _num_chunks_left_rst;
end
endmodule

// BitwiseIntConcat #(UPPER_TO: 2, LOWER_BITS: 2)
module BitwiseIntConcat_UPPER_TO_2_LOWER_BITS_2(
	input clk,
	input wire[0:0] upper,
	input wire[1:0] lower,
	output /*mux_wire*/ logic[2:0] v
);

/*mux_wire*/ logic[2:0] v_bits;
/*mux_wire*/ logic[1:0] _UIntToBits_value;
wire[1:0] _UIntToBits_bits;
/*mux_wire*/ logic[0:0] _UIntToBits_2_value;
wire[0:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[2:0] _FromBits_bits;
wire[2:0] _FromBits_value;
UIntToBits_NUM_BITS_2 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_1 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_8 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 3'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 3'bxxx;
	for(int _v0 = 0; _v0 < 2; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
v_bits[2 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 2'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 1'dx;
	_UIntToBits_2_value = upper;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_UIntToBits_2_value = _UIntToBits_2_value;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 3'bxxx;
	_FromBits_bits = v_bits;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 8))
module FromBits_T_type_int_FROM_0_TO_8(
	input clk,
	input wire[2:0] bits,
	output /*mux_wire*/ logic[2:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 1)
module UIntToBits_NUM_BITS_1(
	input clk,
	input wire[0:0] value,
	output /*mux_wire*/ logic[0:0] bits
);

	assign bits = value;
endmodule

// UIntToBits #(NUM_BITS: 2)
module UIntToBits_NUM_BITS_2(
	input clk,
	input wire[1:0] value,
	output /*mux_wire*/ logic[1:0] bits
);

	assign bits = value;
endmodule

// BitwiseIntSplit #(TO: 65539, LOWER_BITS: 2)
module BitwiseIntSplit_TO_65539_LOWER_BITS_2(
	input clk,
	input wire[16:0] v,
	output /*mux_wire*/ logic[14:0] upper,
	output /*mux_wire*/ logic[1:0] lower
);

genvar _g0;
/*mux_wire*/ logic[16:0] v_bits;
/*mux_wire*/ logic[16:0] _UIntToBits_value;
wire[16:0] _UIntToBits_bits;
wire[1:0] _2;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[1:0] _BitsToUInt_bits;
wire[1:0] _BitsToUInt_value;
wire[14:0] _3;
generate
for(_g0 = 0; _g0 < 15; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[2 + _g0];
end
endgenerate
/*mux_wire*/ logic[14:0] _FromBits_bits;
wire[14:0] _FromBits_value;
UIntToBits_NUM_BITS_17 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_2 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_16385 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 15'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 2'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 17'bxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 17'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 2'bxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 15'bxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 16385))
module FromBits_T_type_int_FROM_0_TO_16385(
	input clk,
	input wire[14:0] bits,
	output /*mux_wire*/ logic[14:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 17)
module UIntToBits_NUM_BITS_17(
	input clk,
	input wire[16:0] value,
	output /*mux_wire*/ logic[16:0] bits
);

	assign bits = value;
endmodule

// BitwiseIntSplit #(TO: 9223372036854775808, LOWER_BITS: 2)
module BitwiseIntSplit_TO_9223372036854775808_LOWER_BITS_2(
	input clk,
	input wire[62:0] v,
	output /*mux_wire*/ logic[60:0] upper,
	output /*mux_wire*/ logic[1:0] lower
);

genvar _g0;
/*mux_wire*/ logic[62:0] v_bits;
/*mux_wire*/ logic[62:0] _UIntToBits_value;
wire[62:0] _UIntToBits_bits;
wire[1:0] _2;
generate
for(_g0 = 0; _g0 < 2; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[1:0] _BitsToUInt_bits;
wire[1:0] _BitsToUInt_value;
wire[60:0] _3;
generate
for(_g0 = 0; _g0 < 61; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[2 + _g0];
end
endgenerate
/*mux_wire*/ logic[60:0] _FromBits_bits;
wire[60:0] _FromBits_value;
UIntToBits_NUM_BITS_63 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_2 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_2305843009213693952 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 61'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 2'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 63'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 63'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 2'bxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 61'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 2305843009213693952))
module FromBits_T_type_int_FROM_0_TO_2305843009213693952(
	input clk,
	input wire[60:0] bits,
	output /*mux_wire*/ logic[60:0] value
);

assign value = bits;
endmodule

// BitsToUInt #(NUM_BITS: 2)
module BitsToUInt_NUM_BITS_2(
	input clk,
	input wire[1:0] bits,
	output /*mux_wire*/ logic[1:0] value
);

	assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 63)
module UIntToBits_NUM_BITS_63(
	input clk,
	input wire[62:0] value,
	output /*mux_wire*/ logic[62:0] bits
);

	assign bits = value;
endmodule

// IntNarrow #(FROM_I: -3, TO_I: 8, FROM: 0, TO: 5)
module IntNarrow_FROM_I_3_TO_I_8_FROM_0_TO_5(
	input clk,
	input wire signed[3:0] in,
	output /*mux_wire*/ logic[2:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: -1, TO_I: 3640, FROM: 0, TO: 3384)
module IntNarrow_FROM_I_1_TO_I_3640_FROM_0_TO_3384(
	input clk,
	input wire signed[12:0] in,
	output /*mux_wire*/ logic[11:0] out
);

	assign out = in;
endmodule

// Ternary #(T: type int #(FROM: 0, TO: 257))
module Ternary_T_type_int_FROM_0_TO_257(
	input clk,
	input wire cond,
	input wire[8:0] a,
	input wire[8:0] b,
	output /*mux_wire*/ logic[8:0] o
);

always_comb begin // combinatorial o
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	o = 9'dx;
	if(cond) o = a;
	if(!cond) o = b;
end
endmodule

// BoolToInt #()
module BoolToInt(
	input clk,
	input wire i,
	output /*mux_wire*/ logic[0:0] o
);

always_comb begin // combinatorial o
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	o = 1'dx;
	if(i) o = 1'd1;
	if(!i) o = 1'd0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	o = o;
end
endmodule

// IntNarrow #(FROM_I: -256, TO_I: 16386, FROM: 0, TO: 16387)
module IntNarrow_FROM_I_256_TO_I_16386_FROM_0_TO_16387(
	input clk,
	input wire signed[15:0] in,
	output /*mux_wire*/ logic[14:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 2305843009213694208, FROM: 0, TO: 2305843009213693952)
module IntNarrow_FROM_I_0_TO_I_2305843009213694208_FROM_0_TO_2305843009213693952(
	input clk,
	input wire[61:0] in,
	output /*mux_wire*/ logic[60:0] out
);

	assign out = in;
endmodule

// BitwiseIntConcat #(UPPER_TO: 9007199254740993, LOWER_BITS: 8)
module BitwiseIntConcat_UPPER_TO_9007199254740993_LOWER_BITS_8(
	input clk,
	input wire[53:0] upper,
	input wire[7:0] lower,
	output /*mux_wire*/ logic[61:0] v
);

/*mux_wire*/ logic[61:0] v_bits;
/*mux_wire*/ logic[7:0] _UIntToBits_value;
wire[7:0] _UIntToBits_bits;
/*mux_wire*/ logic[53:0] _UIntToBits_2_value;
wire[53:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[61:0] _FromBits_bits;
wire[61:0] _FromBits_value;
UIntToBits_NUM_BITS_8 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_54 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_2305843009213694208 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 62'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 62'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 54; _v0 = _v0 + 1) begin
v_bits[8 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 8'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 54'dx;
	_UIntToBits_2_value = upper;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 62'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 2305843009213694208))
module FromBits_T_type_int_FROM_0_TO_2305843009213694208(
	input clk,
	input wire[61:0] bits,
	output /*mux_wire*/ logic[61:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 54)
module UIntToBits_NUM_BITS_54(
	input clk,
	input wire[53:0] value,
	output /*mux_wire*/ logic[53:0] bits
);

	assign bits = value;
endmodule

// UIntToBits #(NUM_BITS: 8)
module UIntToBits_NUM_BITS_8(
	input clk,
	input wire[7:0] value,
	output /*mux_wire*/ logic[7:0] bits
);

	assign bits = value;
endmodule

// LatencyOffset #(T: type bool #(), OFFSET: 384)
module LatencyOffset_T_type_bool_OFFSET_384(
	input clk,
	input wire in,
	output /*mux_wire*/ logic out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 16387, FROM: 1, TO: 257)
module IntNarrow_FROM_I_0_TO_I_16387_FROM_1_TO_257(
	input clk,
	input wire[14:0] in,
	output /*mux_wire*/ logic[8:0] out
);

	assign out = in;
endmodule

// BitwiseIntSplit #(TO: 2305843009213693952, LOWER_BITS: 8)
module BitwiseIntSplit_TO_2305843009213693952_LOWER_BITS_8(
	input clk,
	input wire[60:0] v,
	output /*mux_wire*/ logic[52:0] upper,
	output /*mux_wire*/ logic[7:0] lower
);

genvar _g0;
/*mux_wire*/ logic[60:0] v_bits;
/*mux_wire*/ logic[60:0] _UIntToBits_value;
wire[60:0] _UIntToBits_bits;
wire[7:0] _2;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _2[_g0] = v_bits[_g0];
end
endgenerate
/*mux_wire*/ logic[7:0] _BitsToUInt_bits;
wire[7:0] _BitsToUInt_value;
wire[52:0] _3;
generate
for(_g0 = 0; _g0 < 53; _g0 = _g0 + 1) begin
assign _3[_g0] = v_bits[8 + _g0];
end
endgenerate
/*mux_wire*/ logic[52:0] _FromBits_bits;
wire[52:0] _FromBits_value;
UIntToBits_NUM_BITS_61 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
BitsToUInt_NUM_BITS_8 BitsToUInt(
	.clk(clk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
FromBits_T_type_int_FROM_0_TO_9007199254740992 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial upper
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	upper = 53'dx;
	upper = _FromBits_value;
end
always_comb begin // combinatorial lower
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	lower = 8'dx;
	lower = _BitsToUInt_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 61'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	v_bits = _UIntToBits_bits;
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 61'dx;
	_UIntToBits_value = v;
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 8'bxxxxxxxx;
	_BitsToUInt_bits = _2;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 53'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = _3;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 9007199254740992))
module FromBits_T_type_int_FROM_0_TO_9007199254740992(
	input clk,
	input wire[52:0] bits,
	output /*mux_wire*/ logic[52:0] value
);

assign value = bits;
endmodule

// BitsToUInt #(NUM_BITS: 8)
module BitsToUInt_NUM_BITS_8(
	input clk,
	input wire[7:0] bits,
	output /*mux_wire*/ logic[7:0] value
);

	assign value = bits;
endmodule

// BitwiseIntConcat #(UPPER_TO: 2305843009213693952, LOWER_BITS: 3)
module BitwiseIntConcat_UPPER_TO_2305843009213693952_LOWER_BITS_3(
	input clk,
	input wire[60:0] upper,
	input wire[2:0] lower,
	output /*mux_wire*/ logic[63:0] v
);

/*mux_wire*/ logic[63:0] v_bits;
/*mux_wire*/ logic[2:0] _UIntToBits_value;
wire[2:0] _UIntToBits_bits;
/*mux_wire*/ logic[60:0] _UIntToBits_2_value;
wire[60:0] _UIntToBits_2_bits;
/*mux_wire*/ logic[63:0] _FromBits_bits;
wire[63:0] _FromBits_value;
UIntToBits_NUM_BITS_3 UIntToBits(
	.clk(clk),
	.value(_UIntToBits_value),
	.bits(_UIntToBits_bits)
);
UIntToBits_NUM_BITS_61 UIntToBits_2(
	.clk(clk),
	.value(_UIntToBits_2_value),
	.bits(_UIntToBits_2_bits)
);
FromBits_T_type_int_FROM_0_TO_18446744073709551616 FromBits(
	.clk(clk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v = 64'dx;
	v = _FromBits_value;
end
always_comb begin // combinatorial v_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	v_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 3; _v0 = _v0 + 1) begin
v_bits[_v0] = _UIntToBits_bits[_v0];
end
	for(int _v0 = 0; _v0 < 61; _v0 = _v0 + 1) begin
v_bits[3 + _v0] = _UIntToBits_2_bits[_v0];
end
end
always_comb begin // combinatorial _UIntToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_value = 3'dx;
	_UIntToBits_value = lower;
end
always_comb begin // combinatorial _UIntToBits_2_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_UIntToBits_2_value = 61'dx;
	_UIntToBits_2_value = upper;
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_FromBits_bits = v_bits;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 18446744073709551616))
module FromBits_T_type_int_FROM_0_TO_18446744073709551616(
	input clk,
	input wire[63:0] bits,
	output /*mux_wire*/ logic[63:0] value
);

assign value = bits;
endmodule

// UIntToBits #(NUM_BITS: 61)
module UIntToBits_NUM_BITS_61(
	input clk,
	input wire[60:0] value,
	output /*mux_wire*/ logic[60:0] bits
);

	assign bits = value;
endmodule

// UIntToBits #(NUM_BITS: 3)
module UIntToBits_NUM_BITS_3(
	input clk,
	input wire[2:0] value,
	output /*mux_wire*/ logic[2:0] bits
);

	assign bits = value;
endmodule

// SlowState #(T: type int #(FROM: 0, TO: 16387), RESET_TO: 0, OLD_DELAY: 2, NEW_DELAY: 0)
module SlowState_T_type_int_FROM_0_TO_16387_RESET_TO_0_OLD_DELAY_2_NEW_DELAY_0(
	input clk,
	input wire rst,
	output /*state*/ logic[14:0] old,
	output /*mux_wire*/ logic may_update,
	input wire update,
	input wire[14:0] new_1
);

genvar _g0;
/*mux_wire*/ logic _cross_rst_in;
/*mux_wire*/ logic[14:0] new_s;
/*mux_wire*/ logic update_s;
/*mux_wire*/ logic update_old;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
/*mux_wire*/ logic[14:0] new_old;
/*mux_wire*/ logic[14:0] _LatencyOffset_2_in;
wire[14:0] _LatencyOffset_2_out;
wire _cross_rst_out;
/*latency*/ logic __cross_rst_out_N1; always_ff @(posedge clk) begin __cross_rst_out_N1 <= _cross_rst_out; end
/*latency*/ logic __cross_rst_out_D0; always_ff @(posedge clk) begin __cross_rst_out_D0 <= __cross_rst_out_N1; end
/*state*/ logic[1:0] cooldown;
wire _8 = cooldown[0];
wire _11;
assign _11 = update_s | __cross_rst_out_D0;
/*mux_wire*/ logic _Repeat_v;
wire[1:0] _Repeat_result;
wire[0:0] _12;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _12[_g0] = cooldown[1 + _g0];
end
endgenerate
CrossDomain_T_type_bool cross_rst(
	.in_clk(clk),
	.in(_cross_rst_in),
	.out(_cross_rst_out)
);
LatencyOffset_T_type_bool_OFFSET_2 LatencyOffset(
	.clk(clk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
LatencyOffset_T_type_int_FROM_0_TO_16387_OFFSET_2 LatencyOffset_2(
	.clk(clk),
	.in(_LatencyOffset_2_in),
	.out(_LatencyOffset_2_out)
);
Repeat_T_type_bool_SIZE_2 Repeat(
	.clk(clk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
always_comb begin // combinatorial _cross_rst_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_rst_in = 1'bx;
	_cross_rst_in = rst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_rst_in = _cross_rst_in;
end
always_ff @(posedge clk) begin // state old
	if(_cross_rst_out) old <= 15'd0;
	if(!_cross_rst_out) if(update_old) old <= new_old;
end
always_comb begin // combinatorial new_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_s = 15'dx;
	if(update) new_s = new_1;
end
always_comb begin // combinatorial update_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_s = 1'bx;
	if(update) update_s = 1'b1;
	if(!update) update_s = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_s = update_s;
end
always_comb begin // combinatorial update_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_old = 1'bx;
	update_old = _LatencyOffset_out;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_old = update_old;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = update_s;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial new_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_old = 15'dx;
	new_old = _LatencyOffset_2_out;
end
always_comb begin // combinatorial _LatencyOffset_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_2_in = 15'dx;
	_LatencyOffset_2_in = new_s;
end
always_comb begin // combinatorial may_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_update = 1'bx;
	may_update = _8;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_update = may_update;
end
always_ff @(posedge clk) begin // state cooldown
	if(_11) cooldown <= _Repeat_result;
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(!_11) cooldown[_v0] <= _12[_v0];
end
	if(!_11) cooldown[1] <= 1'b1;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	if(_11) _Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
endmodule

// LatencyOffset #(T: type int #(FROM: 0, TO: 16387), OFFSET: -2)
module LatencyOffset_T_type_int_FROM_0_TO_16387_OFFSET_2(
	input clk,
	input wire[14:0] in,
	output /*mux_wire*/ logic[14:0] out
);

	assign out = in;
endmodule

// SlowState #(T: type int #(FROM: 0, TO: 2305843009213693952), RESET_TO: 0, OLD_DELAY: 1, NEW_DELAY: 1)
module SlowState_T_type_int_FROM_0_TO_2305843009213693952_RESET_TO_0_OLD_DELAY_1_NEW_DELAY_1(
	input clk,
	input wire rst,
	output /*state*/ logic[60:0] old,
	output /*mux_wire*/ logic may_update,
	input wire update,
	input wire[60:0] new_1
);

/*latency*/ logic _update_D1; always_ff @(posedge clk) begin _update_D1 <= update; end
genvar _g0;
/*mux_wire*/ logic _cross_rst_in;
/*mux_wire*/ logic[60:0] new_s;
/*mux_wire*/ logic update_s;
/*mux_wire*/ logic update_old;
/*mux_wire*/ logic _LatencyOffset_in;
wire _LatencyOffset_out;
/*latency*/ logic __LatencyOffset_out_N1; always_ff @(posedge clk) begin __LatencyOffset_out_N1 <= _LatencyOffset_out; end
/*mux_wire*/ logic[60:0] new_old;
/*mux_wire*/ logic[60:0] _LatencyOffset_2_in;
wire[60:0] _LatencyOffset_2_out;
wire _cross_rst_out;
/*latency*/ logic __cross_rst_out_D0; always_ff @(posedge clk) begin __cross_rst_out_D0 <= _cross_rst_out; end
/*state*/ logic[1:0] cooldown;
wire _8 = cooldown[0];
wire _11;
assign _11 = update_s | __cross_rst_out_D0;
/*mux_wire*/ logic _Repeat_v;
wire[1:0] _Repeat_result;
wire[0:0] _12;
generate
for(_g0 = 0; _g0 < 1; _g0 = _g0 + 1) begin
assign _12[_g0] = cooldown[1 + _g0];
end
endgenerate
CrossDomain_T_type_bool cross_rst(
	.in_clk(clk),
	.in(_cross_rst_in),
	.out(_cross_rst_out)
);
LatencyOffset_T_type_bool_OFFSET_2 LatencyOffset(
	.clk(clk),
	.in(_LatencyOffset_in),
	.out(_LatencyOffset_out)
);
LatencyOffset_T_type_int_FROM_0_TO_2305843009213693952_OFFSET_2 LatencyOffset_2(
	.clk(clk),
	.in(_LatencyOffset_2_in),
	.out(_LatencyOffset_2_out)
);
Repeat_T_type_bool_SIZE_2 Repeat(
	.clk(clk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
always_comb begin // combinatorial _cross_rst_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_rst_in = 1'bx;
	_cross_rst_in = rst;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_rst_in = _cross_rst_in;
end
always_ff @(posedge clk) begin // state old
	if(_cross_rst_out) old <= 61'd0;
	if(!_cross_rst_out) if(update_old) old <= new_old;
end
always_comb begin // combinatorial new_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_s = 61'dx;
	if(_update_D1) new_s = new_1;
end
always_comb begin // combinatorial update_s
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_s = 1'bx;
	if(update) update_s = 1'b1;
	if(!update) update_s = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_s = update_s;
end
always_comb begin // combinatorial update_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	update_old = 1'bx;
	update_old = __LatencyOffset_out_N1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	update_old = update_old;
end
always_comb begin // combinatorial _LatencyOffset_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_in = 1'bx;
	_LatencyOffset_in = update_s;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_LatencyOffset_in = _LatencyOffset_in;
end
always_comb begin // combinatorial new_old
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	new_old = 61'dx;
	new_old = _LatencyOffset_2_out;
end
always_comb begin // combinatorial _LatencyOffset_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_LatencyOffset_2_in = 61'dx;
	_LatencyOffset_2_in = new_s;
end
always_comb begin // combinatorial may_update
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	may_update = 1'bx;
	may_update = _8;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	may_update = may_update;
end
always_ff @(posedge clk) begin // state cooldown
	if(_11) cooldown <= _Repeat_result;
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(!_11) cooldown[_v0] <= _12[_v0];
end
	if(!_11) cooldown[1] <= 1'b1;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	if(_11) _Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
endmodule

// Repeat #(T: type bool #(), SIZE: 2)
module Repeat_T_type_bool_SIZE_2(
	input clk,
	input wire v,
	output /*mux_wire*/ logic[1:0] result
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = 2'bxx;
	result[0] = v;
	result[1] = v;
end
endmodule

// LatencyOffset #(T: type int #(FROM: 0, TO: 2305843009213693952), OFFSET: -2)
module LatencyOffset_T_type_int_FROM_0_TO_2305843009213693952_OFFSET_2(
	input clk,
	input wire[60:0] in,
	output /*mux_wire*/ logic[60:0] out
);

	assign out = in;
endmodule

// LatencyOffset #(T: type bool #(), OFFSET: -2)
module LatencyOffset_T_type_bool_OFFSET_2(
	input clk,
	input wire in,
	output /*mux_wire*/ logic out
);

	assign out = in;
endmodule

// combined_axi_ctrl_reader_writer #()
module combined_axi_ctrl_reader_writer(
	input aclk,
	input wire aresetn,
	input wire[11:0] s_axi_control_awaddr,
	input wire s_axi_control_awvalid,
	output /*mux_wire*/ logic s_axi_control_awready,
	input wire[31:0] s_axi_control_wdata,
	input wire[3:0] s_axi_control_wstrb,
	input wire s_axi_control_wvalid,
	output /*mux_wire*/ logic s_axi_control_wready,
	output /*mux_wire*/ logic[1:0] s_axi_control_bresp,
	output /*mux_wire*/ logic s_axi_control_bvalid,
	input wire s_axi_control_bready,
	input wire[11:0] s_axi_control_araddr,
	input wire s_axi_control_arvalid,
	output /*mux_wire*/ logic s_axi_control_arready,
	output /*mux_wire*/ logic[31:0] s_axi_control_rdata,
	output /*mux_wire*/ logic[1:0] s_axi_control_rresp,
	output /*mux_wire*/ logic s_axi_control_rvalid,
	input wire s_axi_control_rready,
	output /*mux_wire*/ logic m_axi_awvalid,
	input wire m_axi_awready,
	output /*mux_wire*/ logic[63:0] m_axi_awaddr,
	output /*mux_wire*/ logic[7:0] m_axi_awlen,
	output /*mux_wire*/ logic[2:0] m_axi_awsize,
	output /*mux_wire*/ logic[1:0] m_axi_awburst,
	output /*mux_wire*/ logic[2:0] m_axi_awprot,
	output /*mux_wire*/ logic[3:0] m_axi_awcache,
	output /*mux_wire*/ logic[3:0] m_axi_awqos,
	output /*mux_wire*/ logic m_axi_awlock,
	output /*mux_wire*/ logic[3:0] m_axi_awregion,
	output /*mux_wire*/ logic m_axi_wvalid,
	input wire m_axi_wready,
	output /*mux_wire*/ logic[31:0] m_axi_wdata,
	output /*mux_wire*/ logic[3:0] m_axi_wstrb,
	output /*mux_wire*/ logic m_axi_wlast,
	input wire m_axi_bvalid,
	output /*mux_wire*/ logic m_axi_bready,
	input wire[1:0] m_axi_bresp,
	output /*mux_wire*/ logic m_axi_arvalid,
	input wire m_axi_arready,
	output /*mux_wire*/ logic[63:0] m_axi_araddr,
	output /*mux_wire*/ logic[7:0] m_axi_arlen,
	output /*mux_wire*/ logic[2:0] m_axi_arsize,
	output /*mux_wire*/ logic[1:0] m_axi_arburst,
	output /*mux_wire*/ logic[2:0] m_axi_arprot,
	output /*mux_wire*/ logic[3:0] m_axi_arcache,
	output /*mux_wire*/ logic[3:0] m_axi_arqos,
	output /*mux_wire*/ logic m_axi_arlock,
	output /*mux_wire*/ logic[3:0] m_axi_arregion,
	input wire m_axi_rvalid,
	output /*mux_wire*/ logic m_axi_rready,
	input wire[31:0] m_axi_rdata,
	input wire[1:0] m_axi_rresp,
	input wire m_axi_rlast
);

/*mux_wire*/ logic _ctrl_aresetn;
wire _ctrl_awready;
wire _ctrl_wready;
wire[1:0] _ctrl_bresp;
wire _ctrl_bvalid;
wire _ctrl_arready;
wire[31:0] _ctrl_rdata;
wire[1:0] _ctrl_rresp;
wire _ctrl_rvalid;
/*mux_wire*/ logic[11:0] _ctrl_awaddr;
/*mux_wire*/ logic _ctrl_awvalid;
/*mux_wire*/ logic[31:0] _ctrl_wdata;
/*mux_wire*/ logic[3:0] _ctrl_wstrb;
/*mux_wire*/ logic _ctrl_wvalid;
/*mux_wire*/ logic _ctrl_bready;
/*mux_wire*/ logic[11:0] _ctrl_araddr;
/*mux_wire*/ logic _ctrl_arvalid;
/*mux_wire*/ logic _ctrl_rready;
/*mux_wire*/ logic _reader_aresetn;
/*mux_wire*/ logic _writer_aresetn;
wire _writer_awvalid;
wire[63:0] _writer_awaddr;
wire[7:0] _writer_awlen;
wire[2:0] _writer_awsize;
wire[1:0] _writer_awburst;
wire[2:0] _writer_awprot;
wire[3:0] _writer_awcache;
wire[3:0] _writer_awqos;
wire _writer_awlock;
wire[3:0] _writer_awregion;
wire _writer_wvalid;
wire[31:0] _writer_wdata;
wire[3:0] _writer_wstrb;
wire _writer_wlast;
wire _writer_bready;
/*mux_wire*/ logic _writer_awready;
/*mux_wire*/ logic _writer_wready;
/*mux_wire*/ logic _writer_bvalid;
/*mux_wire*/ logic[1:0] _writer_bresp;
wire _reader_arvalid;
wire[63:0] _reader_araddr;
wire[7:0] _reader_arlen;
wire[2:0] _reader_arsize;
wire[1:0] _reader_arburst;
wire[2:0] _reader_arprot;
wire[3:0] _reader_arcache;
wire[3:0] _reader_arqos;
wire _reader_arlock;
wire[3:0] _reader_arregion;
wire _reader_rready;
/*mux_wire*/ logic _reader_arready;
/*mux_wire*/ logic _reader_rvalid;
/*mux_wire*/ logic[31:0] _reader_rdata;
/*mux_wire*/ logic[1:0] _reader_rresp;
/*mux_wire*/ logic _reader_rlast;
/*state*/ logic[1:0] addr_state;
/*state*/ logic[2:0] data_state;
/*mux_wire*/ logic[63:0] addr_a_bits;
wire[31:0] _ctrl_input_regs[7:0];
wire[31:0] _56 = _ctrl_input_regs[0];
wire[31:0] _57 = _ctrl_input_regs[1];
/*mux_wire*/ logic[63:0] addr_b_bits;
wire[31:0] _58 = _ctrl_input_regs[2];
wire[31:0] _59 = _ctrl_input_regs[3];
/*mux_wire*/ logic[63:0] addr_c_bits;
wire[31:0] _60 = _ctrl_input_regs[4];
wire[31:0] _61 = _ctrl_input_regs[5];
/*mux_wire*/ logic[63:0] addr_d_bits;
wire[31:0] _62 = _ctrl_input_regs[6];
wire[31:0] _63 = _ctrl_input_regs[7];
wire _65;
assign _65 = addr_state == 1'd1;
/*mux_wire*/ logic[63:0] _BitsToUInt_bits;
wire[63:0] _BitsToUInt_value;
/*mux_wire*/ logic _reader_request;
/*mux_wire*/ logic[63:0] _reader_addr;
wire _reader_fire;
wire _70;
assign _70 = addr_state == 2'd2;
/*mux_wire*/ logic[63:0] _BitsToUInt_2_bits;
wire[63:0] _BitsToUInt_2_value;
/*state*/ logic[31:0] stored_a[7:0];
/*state*/ logic[31:0] stored_b[7:0];
/*mux_wire*/ logic[31:0] c[7:0];
/*mux_wire*/ logic[31:0] d[7:0];
wire[31:0] _73 = stored_a[0];
wire[31:0] _74 = stored_b[0];
wire[32:0] _75;
assign _75 = _73 + _74;
wire[31:0] _76;
assign _76 = _75; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _77 = stored_a[0];
wire[31:0] _78 = stored_b[0];
wire[63:0] _79;
assign _79 = _77 * _78;
wire[31:0] _80;
assign _80 = _79; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _81 = stored_a[1];
wire[31:0] _82 = stored_b[1];
wire[32:0] _83;
assign _83 = _81 + _82;
wire[31:0] _84;
assign _84 = _83; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _85 = stored_a[1];
wire[31:0] _86 = stored_b[1];
wire[63:0] _87;
assign _87 = _85 * _86;
wire[31:0] _88;
assign _88 = _87; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _89 = stored_a[2];
wire[31:0] _90 = stored_b[2];
wire[32:0] _91;
assign _91 = _89 + _90;
wire[31:0] _92;
assign _92 = _91; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _93 = stored_a[2];
wire[31:0] _94 = stored_b[2];
wire[63:0] _95;
assign _95 = _93 * _94;
wire[31:0] _96;
assign _96 = _95; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _97 = stored_a[3];
wire[31:0] _98 = stored_b[3];
wire[32:0] _99;
assign _99 = _97 + _98;
wire[31:0] _100;
assign _100 = _99; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _101 = stored_a[3];
wire[31:0] _102 = stored_b[3];
wire[63:0] _103;
assign _103 = _101 * _102;
wire[31:0] _104;
assign _104 = _103; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _105 = stored_a[4];
wire[31:0] _106 = stored_b[4];
wire[32:0] _107;
assign _107 = _105 + _106;
wire[31:0] _108;
assign _108 = _107; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _109 = stored_a[4];
wire[31:0] _110 = stored_b[4];
wire[63:0] _111;
assign _111 = _109 * _110;
wire[31:0] _112;
assign _112 = _111; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _113 = stored_a[5];
wire[31:0] _114 = stored_b[5];
wire[32:0] _115;
assign _115 = _113 + _114;
wire[31:0] _116;
assign _116 = _115; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _117 = stored_a[5];
wire[31:0] _118 = stored_b[5];
wire[63:0] _119;
assign _119 = _117 * _118;
wire[31:0] _120;
assign _120 = _119; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _121 = stored_a[6];
wire[31:0] _122 = stored_b[6];
wire[32:0] _123;
assign _123 = _121 + _122;
wire[31:0] _124;
assign _124 = _123; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _125 = stored_a[6];
wire[31:0] _126 = stored_b[6];
wire[63:0] _127;
assign _127 = _125 * _126;
wire[31:0] _128;
assign _128 = _127; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _129 = stored_a[7];
wire[31:0] _130 = stored_b[7];
wire[32:0] _131;
assign _131 = _129 + _130;
wire[31:0] _132;
assign _132 = _131; // == mod 4294967296 (target is 32 bits wide)
wire[31:0] _133 = stored_a[7];
wire[31:0] _134 = stored_b[7];
wire[63:0] _135;
assign _135 = _133 * _134;
wire[31:0] _136;
assign _136 = _135; // == mod 4294967296 (target is 32 bits wide)
wire _138;
assign _138 = data_state == 1'd1;
/*mux_wire*/ logic success;
/*mux_wire*/ logic[31:0] data[7:0];
/*mux_wire*/ logic _reader_read;
wire _reader_read_valid;
wire[31:0] _reader_data[7:0];
wire _144;
assign _144 = data_state == 2'd2;
/*mux_wire*/ logic success_2;
/*mux_wire*/ logic[31:0] data_2[7:0];
wire _149;
assign _149 = data_state == 2'd3;
/*mux_wire*/ logic[63:0] _BitsToUInt_3_bits;
wire[63:0] _BitsToUInt_3_value;
/*mux_wire*/ logic _writer_write;
/*mux_wire*/ logic[63:0] _writer_addr;
/*mux_wire*/ logic[31:0] _writer_data[7:0];
wire _writer_write_success;
wire _155;
assign _155 = data_state == 3'd4;
/*mux_wire*/ logic[63:0] _BitsToUInt_4_bits;
wire[63:0] _BitsToUInt_4_value;
wire _160;
assign _160 = data_state == 3'd5;
wire _writer_has_outstanding_writes;
wire _162;
assign _162 = !_writer_has_outstanding_writes;
/*mux_wire*/ logic _ctrl_finish;
/*mux_wire*/ logic[31:0] _ctrl_output_regs[0:0];
localparam[31:0] _165[0:0] = '{32'b11011110101011011011111011101111};
wire _ctrl_start;
wire _167;
assign _167 = !aresetn;
axi_ctrl_slave_NUM_INPUT_REGS_8_NUM_OUTPUT_REGS_1_ADDR_WIDTH_12_AXI_WIDTH_32 ctrl(
	.aclk(aclk),
	.aresetn(_ctrl_aresetn),
	.awaddr(_ctrl_awaddr),
	.awvalid(_ctrl_awvalid),
	.awready(_ctrl_awready),
	.wdata(_ctrl_wdata),
	.wstrb(_ctrl_wstrb),
	.wvalid(_ctrl_wvalid),
	.wready(_ctrl_wready),
	.bresp(_ctrl_bresp),
	.bvalid(_ctrl_bvalid),
	.bready(_ctrl_bready),
	.araddr(_ctrl_araddr),
	.arvalid(_ctrl_arvalid),
	.arready(_ctrl_arready),
	.rdata(_ctrl_rdata),
	.rresp(_ctrl_rresp),
	.rvalid(_ctrl_rvalid),
	.rready(_ctrl_rready),
	.input_regs(_ctrl_input_regs),
	.start(_ctrl_start),
	.finish(_ctrl_finish),
	.output_regs(_ctrl_output_regs)
);
axi_memory_reader_T_type_int_FROM_0_TO_4294967296_8_AXI_WIDTH_32 reader(
	.aclk(aclk),
	.aresetn(_reader_aresetn),
	.arvalid(_reader_arvalid),
	.arready(_reader_arready),
	.araddr(_reader_araddr),
	.arlen(_reader_arlen),
	.arsize(_reader_arsize),
	.arburst(_reader_arburst),
	.arprot(_reader_arprot),
	.arcache(_reader_arcache),
	.arqos(_reader_arqos),
	.arlock(_reader_arlock),
	.arregion(_reader_arregion),
	.rvalid(_reader_rvalid),
	.rready(_reader_rready),
	.rdata(_reader_rdata),
	.rresp(_reader_rresp),
	.rlast(_reader_rlast),
	.request(_reader_request),
	.addr(_reader_addr),
	.fire(_reader_fire),
	.read(_reader_read),
	.read_valid(_reader_read_valid),
	.data(_reader_data)
);
axi_memory_writer_T_type_int_FROM_0_TO_4294967296_8_AXI_WIDTH_32 writer(
	.aclk(aclk),
	.aresetn(_writer_aresetn),
	.awvalid(_writer_awvalid),
	.awready(_writer_awready),
	.awaddr(_writer_awaddr),
	.awlen(_writer_awlen),
	.awsize(_writer_awsize),
	.awburst(_writer_awburst),
	.awprot(_writer_awprot),
	.awcache(_writer_awcache),
	.awqos(_writer_awqos),
	.awlock(_writer_awlock),
	.awregion(_writer_awregion),
	.wvalid(_writer_wvalid),
	.wready(_writer_wready),
	.wdata(_writer_wdata),
	.wstrb(_writer_wstrb),
	.wlast(_writer_wlast),
	.bvalid(_writer_bvalid),
	.bready(_writer_bready),
	.bresp(_writer_bresp),
	.has_outstanding_writes(_writer_has_outstanding_writes),
	.write(_writer_write),
	.addr(_writer_addr),
	.data(_writer_data),
	.write_success(_writer_write_success)
);
BitsToUInt_NUM_BITS_64 BitsToUInt(
	.clk(aclk),
	.bits(_BitsToUInt_bits),
	.value(_BitsToUInt_value)
);
BitsToUInt_NUM_BITS_64 BitsToUInt_2(
	.clk(aclk),
	.bits(_BitsToUInt_2_bits),
	.value(_BitsToUInt_2_value)
);
BitsToUInt_NUM_BITS_64 BitsToUInt_3(
	.clk(aclk),
	.bits(_BitsToUInt_3_bits),
	.value(_BitsToUInt_3_value)
);
BitsToUInt_NUM_BITS_64 BitsToUInt_4(
	.clk(aclk),
	.bits(_BitsToUInt_4_bits),
	.value(_BitsToUInt_4_value)
);
always_comb begin // combinatorial _ctrl_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_aresetn = 1'bx;
	_ctrl_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_aresetn = _ctrl_aresetn;
end
always_comb begin // combinatorial s_axi_control_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_awready = 1'bx;
	s_axi_control_awready = _ctrl_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_awready = s_axi_control_awready;
end
always_comb begin // combinatorial s_axi_control_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_wready = 1'bx;
	s_axi_control_wready = _ctrl_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_wready = s_axi_control_wready;
end
always_comb begin // combinatorial s_axi_control_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bresp = 2'bxx;
	s_axi_control_bresp = _ctrl_bresp;
end
always_comb begin // combinatorial s_axi_control_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_bvalid = 1'bx;
	s_axi_control_bvalid = _ctrl_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_bvalid = s_axi_control_bvalid;
end
always_comb begin // combinatorial s_axi_control_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_arready = 1'bx;
	s_axi_control_arready = _ctrl_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_arready = s_axi_control_arready;
end
always_comb begin // combinatorial s_axi_control_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	s_axi_control_rdata = _ctrl_rdata;
end
always_comb begin // combinatorial s_axi_control_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rresp = 2'bxx;
	s_axi_control_rresp = _ctrl_rresp;
end
always_comb begin // combinatorial s_axi_control_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	s_axi_control_rvalid = 1'bx;
	s_axi_control_rvalid = _ctrl_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	s_axi_control_rvalid = s_axi_control_rvalid;
end
always_comb begin // combinatorial _ctrl_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awaddr = 12'dx;
	_ctrl_awaddr = s_axi_control_awaddr;
end
always_comb begin // combinatorial _ctrl_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_awvalid = 1'bx;
	_ctrl_awvalid = s_axi_control_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_awvalid = _ctrl_awvalid;
end
always_comb begin // combinatorial _ctrl_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_ctrl_wdata = s_axi_control_wdata;
end
always_comb begin // combinatorial _ctrl_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wstrb = 4'bxxxx;
	_ctrl_wstrb = s_axi_control_wstrb;
end
always_comb begin // combinatorial _ctrl_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_wvalid = 1'bx;
	_ctrl_wvalid = s_axi_control_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_wvalid = _ctrl_wvalid;
end
always_comb begin // combinatorial _ctrl_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_bready = 1'bx;
	_ctrl_bready = s_axi_control_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_bready = _ctrl_bready;
end
always_comb begin // combinatorial _ctrl_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_araddr = 12'dx;
	_ctrl_araddr = s_axi_control_araddr;
end
always_comb begin // combinatorial _ctrl_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_arvalid = 1'bx;
	_ctrl_arvalid = s_axi_control_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_arvalid = _ctrl_arvalid;
end
always_comb begin // combinatorial _ctrl_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_rready = 1'bx;
	_ctrl_rready = s_axi_control_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_rready = _ctrl_rready;
end
always_comb begin // combinatorial _reader_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_aresetn = 1'bx;
	_reader_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_aresetn = _reader_aresetn;
end
always_comb begin // combinatorial _writer_aresetn
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_aresetn = 1'bx;
	_writer_aresetn = aresetn;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_aresetn = _writer_aresetn;
end
always_comb begin // combinatorial m_axi_awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awvalid = 1'bx;
	m_axi_awvalid = _writer_awvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_awvalid = m_axi_awvalid;
end
always_comb begin // combinatorial m_axi_awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awaddr = 64'dx;
	m_axi_awaddr = _writer_awaddr;
end
always_comb begin // combinatorial m_axi_awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awlen = 8'dx;
	m_axi_awlen = _writer_awlen;
end
always_comb begin // combinatorial m_axi_awsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awsize = 3'dx;
	m_axi_awsize = _writer_awsize;
end
always_comb begin // combinatorial m_axi_awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awburst = 2'bxx;
	m_axi_awburst = _writer_awburst;
end
always_comb begin // combinatorial m_axi_awprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awprot = 3'bxxx;
	m_axi_awprot = _writer_awprot;
end
always_comb begin // combinatorial m_axi_awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awcache = 4'bxxxx;
	m_axi_awcache = _writer_awcache;
end
always_comb begin // combinatorial m_axi_awqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awqos = 4'dx;
	m_axi_awqos = _writer_awqos;
end
always_comb begin // combinatorial m_axi_awlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awlock = 1'bx;
	m_axi_awlock = _writer_awlock;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_awlock = m_axi_awlock;
end
always_comb begin // combinatorial m_axi_awregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_awregion = 4'dx;
	m_axi_awregion = _writer_awregion;
end
always_comb begin // combinatorial m_axi_wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wvalid = 1'bx;
	m_axi_wvalid = _writer_wvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wvalid = m_axi_wvalid;
end
always_comb begin // combinatorial m_axi_wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	m_axi_wdata = _writer_wdata;
end
always_comb begin // combinatorial m_axi_wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wstrb = 4'bxxxx;
	m_axi_wstrb = _writer_wstrb;
end
always_comb begin // combinatorial m_axi_wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_wlast = 1'bx;
	m_axi_wlast = _writer_wlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_wlast = m_axi_wlast;
end
always_comb begin // combinatorial m_axi_bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_bready = 1'bx;
	m_axi_bready = _writer_bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_bready = m_axi_bready;
end
always_comb begin // combinatorial _writer_awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_awready = 1'bx;
	_writer_awready = m_axi_awready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_awready = _writer_awready;
end
always_comb begin // combinatorial _writer_wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_wready = 1'bx;
	_writer_wready = m_axi_wready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_wready = _writer_wready;
end
always_comb begin // combinatorial _writer_bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bvalid = 1'bx;
	_writer_bvalid = m_axi_bvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_bvalid = _writer_bvalid;
end
always_comb begin // combinatorial _writer_bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_bresp = 2'bxx;
	_writer_bresp = m_axi_bresp;
end
always_comb begin // combinatorial m_axi_arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arvalid = 1'bx;
	m_axi_arvalid = _reader_arvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arvalid = m_axi_arvalid;
end
always_comb begin // combinatorial m_axi_araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_araddr = 64'dx;
	m_axi_araddr = _reader_araddr;
end
always_comb begin // combinatorial m_axi_arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlen = 8'dx;
	m_axi_arlen = _reader_arlen;
end
always_comb begin // combinatorial m_axi_arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arsize = 3'dx;
	m_axi_arsize = _reader_arsize;
end
always_comb begin // combinatorial m_axi_arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arburst = 2'bxx;
	m_axi_arburst = _reader_arburst;
end
always_comb begin // combinatorial m_axi_arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arprot = 3'bxxx;
	m_axi_arprot = _reader_arprot;
end
always_comb begin // combinatorial m_axi_arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arcache = 4'bxxxx;
	m_axi_arcache = _reader_arcache;
end
always_comb begin // combinatorial m_axi_arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arqos = 4'dx;
	m_axi_arqos = _reader_arqos;
end
always_comb begin // combinatorial m_axi_arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arlock = 1'bx;
	m_axi_arlock = _reader_arlock;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_arlock = m_axi_arlock;
end
always_comb begin // combinatorial m_axi_arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_arregion = 4'dx;
	m_axi_arregion = _reader_arregion;
end
always_comb begin // combinatorial m_axi_rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	m_axi_rready = 1'bx;
	m_axi_rready = _reader_rready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	m_axi_rready = m_axi_rready;
end
always_comb begin // combinatorial _reader_arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_arready = 1'bx;
	_reader_arready = m_axi_arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_arready = _reader_arready;
end
always_comb begin // combinatorial _reader_rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rvalid = 1'bx;
	_reader_rvalid = m_axi_rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rvalid = _reader_rvalid;
end
always_comb begin // combinatorial _reader_rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	_reader_rdata = m_axi_rdata;
end
always_comb begin // combinatorial _reader_rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rresp = 2'bxx;
	_reader_rresp = m_axi_rresp;
end
always_comb begin // combinatorial _reader_rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_rlast = 1'bx;
	_reader_rlast = m_axi_rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_rlast = _reader_rlast;
end
always_ff @(posedge aclk) begin // state addr_state
	if(_65) if(_reader_fire) addr_state <= 2'd2;
	if(!_65) if(_70) if(_reader_fire) addr_state <= 1'd0;
	if(_ctrl_start) addr_state <= 1'd1;
	if(_167) addr_state <= 1'd0;
end
always_ff @(posedge aclk) begin // state data_state
	if(_138) if(success) data_state <= 2'd2;
	if(!_138) if(_144) if(success_2) data_state <= 2'd3;
	if(!_138) if(!_144) if(_149) if(_writer_write_success) data_state <= 3'd4;
	if(!_138) if(!_144) if(!_149) if(_155) if(_writer_write_success) data_state <= 3'd5;
	if(!_138) if(!_144) if(!_149) if(!_155) if(_160) if(_162) data_state <= 1'd0;
	if(_ctrl_start) data_state <= 1'd1;
	if(_167) data_state <= 1'd0;
end
always_comb begin // combinatorial addr_a_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	addr_a_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[_v0] = _56[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_a_bits[32 + _v0] = _57[_v0];
end
end
always_comb begin // combinatorial addr_b_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	addr_b_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_b_bits[_v0] = _58[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_b_bits[32 + _v0] = _59[_v0];
end
end
always_comb begin // combinatorial addr_c_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	addr_c_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_c_bits[_v0] = _60[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_c_bits[32 + _v0] = _61[_v0];
end
end
always_comb begin // combinatorial addr_d_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	addr_d_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_d_bits[_v0] = _62[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
addr_d_bits[32 + _v0] = _63[_v0];
end
end
always_comb begin // combinatorial _BitsToUInt_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_65) _BitsToUInt_bits = addr_a_bits;
end
always_comb begin // combinatorial _reader_request
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_request = 1'bx;
	_reader_request = 1'b0;
	if(_65) _reader_request = 1'b1;
	if(!_65) if(_70) _reader_request = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_request = _reader_request;
end
always_comb begin // combinatorial _reader_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_addr = 64'dx;
	if(_65) _reader_addr = _BitsToUInt_value;
	if(!_65) if(_70) _reader_addr = _BitsToUInt_2_value;
end
always_comb begin // combinatorial _BitsToUInt_2_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_2_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(!_65) if(_70) _BitsToUInt_2_bits = addr_b_bits;
end
always_ff @(posedge aclk) begin // state stored_a
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_138) if(success) stored_a[_v0] <= data[_v0];
end
end
always_ff @(posedge aclk) begin // state stored_b
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(!_138) if(_144) if(success_2) stored_b[_v0] <= data_2[_v0];
end
end
always_comb begin // combinatorial c
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	c = '{32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx};
	c[0] = _76;
	c[1] = _84;
	c[2] = _92;
	c[3] = _100;
	c[4] = _108;
	c[5] = _116;
	c[6] = _124;
	c[7] = _132;
end
always_comb begin // combinatorial d
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	d = '{32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx};
	d[0] = _80;
	d[1] = _88;
	d[2] = _96;
	d[3] = _104;
	d[4] = _112;
	d[5] = _120;
	d[6] = _128;
	d[7] = _136;
end
always_comb begin // combinatorial success
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	success = 1'bx;
	if(_138) success = _reader_read_valid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	success = success;
end
always_comb begin // combinatorial data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	data = '{32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_138) data[_v0] = _reader_data[_v0];
end
end
always_comb begin // combinatorial _reader_read
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_reader_read = 1'bx;
	_reader_read = 1'b0;
	if(_138) _reader_read = 1'b1;
	if(!_138) if(_144) _reader_read = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_reader_read = _reader_read;
end
always_comb begin // combinatorial success_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	success_2 = 1'bx;
	if(!_138) if(_144) success_2 = _reader_read_valid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	success_2 = success_2;
end
always_comb begin // combinatorial data_2
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	data_2 = '{32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(!_138) if(_144) data_2[_v0] = _reader_data[_v0];
end
end
always_comb begin // combinatorial _BitsToUInt_3_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_3_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(!_138) if(!_144) if(_149) _BitsToUInt_3_bits = addr_c_bits;
end
always_comb begin // combinatorial _writer_write
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_write = 1'bx;
	_writer_write = 1'b0;
	if(!_138) if(!_144) if(_149) _writer_write = 1'b1;
	if(!_138) if(!_144) if(!_149) if(_155) _writer_write = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_writer_write = _writer_write;
end
always_comb begin // combinatorial _writer_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_addr = 64'dx;
	if(!_138) if(!_144) if(_149) _writer_addr = _BitsToUInt_3_value;
	if(!_138) if(!_144) if(!_149) if(_155) _writer_addr = _BitsToUInt_4_value;
end
always_comb begin // combinatorial _writer_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_writer_data = '{32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(!_138) if(!_144) if(_149) _writer_data[_v0] = c[_v0];
end
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(!_138) if(!_144) if(!_149) if(_155) _writer_data[_v0] = d[_v0];
end
end
always_comb begin // combinatorial _BitsToUInt_4_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_BitsToUInt_4_bits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(!_138) if(!_144) if(!_149) if(_155) _BitsToUInt_4_bits = addr_d_bits;
end
always_comb begin // combinatorial _ctrl_finish
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_finish = 1'bx;
	_ctrl_finish = 1'b0;
	if(!_138) if(!_144) if(!_149) if(!_155) if(_160) if(_162) _ctrl_finish = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_ctrl_finish = _ctrl_finish;
end
always_comb begin // combinatorial _ctrl_output_regs
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ctrl_output_regs = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(!_138) if(!_144) if(!_149) if(!_155) if(_160) if(_162) _ctrl_output_regs[_v0] = _165[_v0];
end
end
endmodule

// BitsToUInt #(NUM_BITS: 64)
module BitsToUInt_NUM_BITS_64(
	input clk,
	input wire[63:0] bits,
	output /*mux_wire*/ logic[63:0] value
);

	assign value = bits;
endmodule

// axi_memory_writer #(T: type int #(FROM: 0, TO: 4294967296)[8], AXI_WIDTH: 32)
module axi_memory_writer_T_type_int_FROM_0_TO_4294967296_8_AXI_WIDTH_32(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic awvalid,
	input wire awready,
	output /*mux_wire*/ logic[63:0] awaddr,
	output /*mux_wire*/ logic[7:0] awlen,
	output /*mux_wire*/ logic[2:0] awsize,
	output /*mux_wire*/ logic[1:0] awburst,
	output /*mux_wire*/ logic[2:0] awprot,
	output /*mux_wire*/ logic[3:0] awcache,
	output /*mux_wire*/ logic[3:0] awqos,
	output /*mux_wire*/ logic awlock,
	output /*mux_wire*/ logic[3:0] awregion,
	output /*mux_wire*/ logic wvalid,
	input wire wready,
	output /*mux_wire*/ logic[31:0] wdata,
	output /*mux_wire*/ logic[3:0] wstrb,
	output /*mux_wire*/ logic wlast,
	input wire bvalid,
	output /*mux_wire*/ logic bready,
	input wire[1:0] bresp,
	output /*mux_wire*/ logic has_outstanding_writes,
	input wire write,
	input wire[63:0] addr,
	input wire[31:0] data[7:0],
	output /*mux_wire*/ logic write_success
);

genvar _g0;
localparam[2:0] _1 = 3'b000;
localparam[3:0] _2 = 4'b0010;
/*mux_wire*/ logic[1:0] _bresp;
/*state*/ logic[255:0] writing_data;
/*state*/ logic writing_data_valid;
/*state*/ logic[7:0] num_outstanding_writes;
wire _9;
assign _9 = num_outstanding_writes != 1'd0;
/*state*/ logic[2:0] cur_data_chunk;
/*mux_wire*/ logic[31:0] parts[7:0];
wire[31:0] _10;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _10[_g0] = writing_data[_g0];
end
endgenerate
wire[31:0] _11;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _11[_g0] = writing_data[32 + _g0];
end
endgenerate
wire[31:0] _12;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _12[_g0] = writing_data[64 + _g0];
end
endgenerate
wire[31:0] _13;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _13[_g0] = writing_data[96 + _g0];
end
endgenerate
wire[31:0] _14;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _14[_g0] = writing_data[128 + _g0];
end
endgenerate
wire[31:0] _15;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _15[_g0] = writing_data[160 + _g0];
end
endgenerate
wire[31:0] _16;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _16[_g0] = writing_data[192 + _g0];
end
endgenerate
wire[31:0] _17;
generate
for(_g0 = 0; _g0 < 32; _g0 = _g0 + 1) begin
assign _17[_g0] = writing_data[224 + _g0];
end
endgenerate
wire[31:0] _19 = parts[cur_data_chunk];
/*mux_wire*/ logic _Repeat_v;
wire[3:0] _Repeat_result;
wire _22;
assign _22 = cur_data_chunk < 3'd7;
wire _23;
assign _23 = !_22;
wire _26;
assign _26 = wvalid & wready;
wire _28;
assign _28 = !wlast;
wire[3:0] _31;
assign _31 = cur_data_chunk + 1'd1;
/*mux_wire*/ logic[3:0] _IntNarrow_in;
wire[2:0] _IntNarrow_out;
wire _34;
assign _34 = awvalid & awready;
localparam[1:0] _38 = 2'b01;
wire _41;
assign _41 = !writing_data_valid;
wire _44;
assign _44 = num_outstanding_writes < 8'd255;
wire _45;
assign _45 = _41 & _44;
wire _48;
assign _48 = awvalid & awready;
wire _51;
assign _51 = awvalid & awready;
/*mux_wire*/ logic[31:0] _ToBits_value[7:0];
wire[255:0] _ToBits_bits;
wire _55;
assign _55 = awvalid & awready;
wire _58;
assign _58 = bvalid & bready;
wire _59;
assign _59 = !_58;
wire _60;
assign _60 = _55 & _59;
/*mux_wire*/ logic[7:0] _IntNarrow_2_in;
wire[7:0] _IntNarrow_2_out;
wire[7:0] _63;
assign _63 = _IntNarrow_2_out + 1'd1;
wire _66;
assign _66 = bvalid & bready;
wire _69;
assign _69 = awvalid & awready;
wire _70;
assign _70 = !_69;
wire _71;
assign _71 = _66 & _70;
/*mux_wire*/ logic[7:0] _IntNarrow_3_in;
wire[7:0] _IntNarrow_3_out;
wire[7:0] _74;
assign _74 = _IntNarrow_3_out - 1'd1;
wire _76;
assign _76 = !aresetn;
Repeat_T_type_bool_SIZE_4 Repeat(
	.clk(aclk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
IntNarrow_FROM_I_1_TO_I_9_FROM_0_TO_7 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
ToBits_T_type_int_FROM_0_TO_4294967296_8 ToBits(
	.clk(aclk),
	.value(_ToBits_value),
	.bits(_ToBits_bits)
);
IntNarrow_FROM_I_0_TO_I_256_FROM_0_TO_255 IntNarrow_2(
	.clk(aclk),
	.in(_IntNarrow_2_in),
	.out(_IntNarrow_2_out)
);
IntNarrow_FROM_I_0_TO_I_256_FROM_1_TO_256 IntNarrow_3(
	.clk(aclk),
	.in(_IntNarrow_3_in),
	.out(_IntNarrow_3_out)
);
always_comb begin // combinatorial awvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awvalid = 1'bx;
	if(write) awvalid = _45;
	if(!write) awvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awvalid = awvalid;
end
always_comb begin // combinatorial awaddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awaddr = 64'dx;
	if(write) awaddr = addr;
end
always_comb begin // combinatorial awlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlen = 8'dx;
	if(write) awlen = 3'd7;
end
always_comb begin // combinatorial awsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awsize = 3'dx;
	awsize = 2'd2;
end
always_comb begin // combinatorial awburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awburst = 2'bxx;
	if(write) awburst = _38;
end
always_comb begin // combinatorial awprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awprot = 3'bxxx;
	awprot = _1;
end
always_comb begin // combinatorial awcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awcache = 4'bxxxx;
	awcache = _2;
end
always_comb begin // combinatorial awqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awqos = 4'dx;
	awqos = 1'd0;
end
always_comb begin // combinatorial awlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awlock = 1'bx;
	awlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awlock = awlock;
end
always_comb begin // combinatorial awregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awregion = 4'dx;
	awregion = 1'd0;
end
always_comb begin // combinatorial wvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wvalid = 1'bx;
	wvalid = writing_data_valid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wvalid = wvalid;
end
always_comb begin // combinatorial wdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	wdata = _19;
end
always_comb begin // combinatorial wstrb
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wstrb = 4'bxxxx;
	wstrb = _Repeat_result;
end
always_comb begin // combinatorial wlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wlast = 1'bx;
	wlast = _23;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wlast = wlast;
end
always_comb begin // combinatorial bready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	bready = 1'bx;
	bready = _9;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	bready = bready;
end
always_comb begin // combinatorial _bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_bresp = 2'bxx;
	_bresp = bresp;
end
always_ff @(posedge aclk) begin // state writing_data
	if(write) if(_51) writing_data <= _ToBits_bits;
end
always_ff @(posedge aclk) begin // state writing_data_valid
	if(_26) if(!_28) writing_data_valid <= 1'b0;
	if(write) if(_51) writing_data_valid <= 1'b1;
	if(_76) writing_data_valid <= 1'b0;
end
always_ff @(posedge aclk) begin // state num_outstanding_writes
	if(_60) num_outstanding_writes <= _63;
	if(!_60) if(_71) num_outstanding_writes <= _74;
	if(_76) num_outstanding_writes <= 1'd0;
end
always_ff @(posedge aclk) begin // state cur_data_chunk
	if(_26) if(_28) cur_data_chunk <= _IntNarrow_out;
	if(_34) cur_data_chunk <= 1'd0;
end
always_comb begin // combinatorial parts
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	parts = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	parts[0] = _10;
	parts[1] = _11;
	parts[2] = _12;
	parts[3] = _13;
	parts[4] = _14;
	parts[5] = _15;
	parts[6] = _16;
	parts[7] = _17;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	_Repeat_v = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 4'dx;
	if(_26) if(_28) _IntNarrow_in = _31;
end
always_comb begin // combinatorial has_outstanding_writes
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	has_outstanding_writes = 1'bx;
	has_outstanding_writes = bready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	has_outstanding_writes = has_outstanding_writes;
end
always_comb begin // combinatorial write_success
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	write_success = 1'bx;
	if(write) write_success = _48;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	write_success = write_success;
end
always_comb begin // combinatorial _ToBits_value
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_ToBits_value = '{32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(write) if(_51) _ToBits_value[_v0] = data[_v0];
end
end
always_comb begin // combinatorial _IntNarrow_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_2_in = 8'dx;
	if(_60) _IntNarrow_2_in = num_outstanding_writes;
end
always_comb begin // combinatorial _IntNarrow_3_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_3_in = 8'dx;
	if(!_60) if(_71) _IntNarrow_3_in = num_outstanding_writes;
end
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 256, FROM: 1, TO: 256)
module IntNarrow_FROM_I_0_TO_I_256_FROM_1_TO_256(
	input clk,
	input wire[7:0] in,
	output /*mux_wire*/ logic[7:0] out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 256, FROM: 0, TO: 255)
module IntNarrow_FROM_I_0_TO_I_256_FROM_0_TO_255(
	input clk,
	input wire[7:0] in,
	output /*mux_wire*/ logic[7:0] out
);

	assign out = in;
endmodule

// ToBits #(T: type int #(FROM: 0, TO: 4294967296)[8])
module ToBits_T_type_int_FROM_0_TO_4294967296_8(
	input clk,
	input wire[31:0] value[7:0],
	output /*mux_wire*/ logic[255:0] bits
);

genvar _g0;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign bits[(_g0) * 32 +: 32] = value[_g0];
end
endgenerate
endmodule

// IntNarrow #(FROM_I: 1, TO_I: 9, FROM: 0, TO: 7)
module IntNarrow_FROM_I_1_TO_I_9_FROM_0_TO_7(
	input clk,
	input wire[3:0] in,
	output /*mux_wire*/ logic[2:0] out
);

	assign out = in;
endmodule

// Repeat #(T: type bool #(), SIZE: 4)
module Repeat_T_type_bool_SIZE_4(
	input clk,
	input wire v,
	output /*mux_wire*/ logic[3:0] result
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = 4'bxxxx;
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
end
endmodule

// axi_memory_reader #(T: type int #(FROM: 0, TO: 4294967296)[8], AXI_WIDTH: 32)
module axi_memory_reader_T_type_int_FROM_0_TO_4294967296_8_AXI_WIDTH_32(
	input aclk,
	input wire aresetn,
	output /*mux_wire*/ logic arvalid,
	input wire arready,
	output /*mux_wire*/ logic[63:0] araddr,
	output /*mux_wire*/ logic[7:0] arlen,
	output /*mux_wire*/ logic[2:0] arsize,
	output /*mux_wire*/ logic[1:0] arburst,
	output /*mux_wire*/ logic[2:0] arprot,
	output /*mux_wire*/ logic[3:0] arcache,
	output /*mux_wire*/ logic[3:0] arqos,
	output /*mux_wire*/ logic arlock,
	output /*mux_wire*/ logic[3:0] arregion,
	input wire rvalid,
	output /*mux_wire*/ logic rready,
	input wire[31:0] rdata,
	input wire[1:0] rresp,
	input wire rlast,
	input wire request,
	input wire[63:0] addr,
	output /*mux_wire*/ logic fire,
	input wire read,
	output /*mux_wire*/ logic read_valid,
	output /*mux_wire*/ logic[31:0] data[7:0]
);

localparam[1:0] _1 = 2'b01;
localparam[2:0] _2 = 3'b000;
localparam[3:0] _3 = 4'b0010;
/*mux_wire*/ logic[1:0] _rresp;
/*mux_wire*/ logic _rlast;
/*mux_wire*/ logic do_read;
/*mux_wire*/ logic do_read_was_valid;
/*mux_wire*/ logic[255:0] do_read_data;
/*state*/ logic[2:0] stored_part_idx;
/*state*/ logic[31:0] stored_parts[6:0];
wire _13;
assign _13 = stored_part_idx < 3'd7;
/*mux_wire*/ logic[2:0] idx;
/*mux_wire*/ logic[2:0] _IntNarrow_in;
wire[2:0] _IntNarrow_out;
wire[2:0] _20;
assign _20 = idx + 1'd1;
wire _25;
assign _25 = rready & rvalid;
wire[31:0] _27 = stored_parts[0];
wire[31:0] _28 = stored_parts[1];
wire[31:0] _29 = stored_parts[2];
wire[31:0] _30 = stored_parts[3];
wire[31:0] _31 = stored_parts[4];
wire[31:0] _32 = stored_parts[5];
wire[31:0] _33 = stored_parts[6];
wire _36;
assign _36 = !aresetn;
/*mux_wire*/ logic[255:0] _FromBits_bits;
wire[31:0] _FromBits_value[7:0];
IntNarrow_FROM_I_0_TO_I_8_FROM_0_TO_7 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
FromBits_T_type_int_FROM_0_TO_4294967296_8 FromBits(
	.clk(aclk),
	.bits(_FromBits_bits),
	.value(_FromBits_value)
);
always_comb begin // combinatorial arvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arvalid = 1'bx;
	if(request) arvalid = 1'b1;
	if(!request) arvalid = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arvalid = arvalid;
end
always_comb begin // combinatorial araddr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	araddr = 64'dx;
	if(request) araddr = addr;
end
always_comb begin // combinatorial arlen
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlen = 8'dx;
	if(request) arlen = 3'd7;
end
always_comb begin // combinatorial arsize
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arsize = 3'dx;
	arsize = 2'd2;
end
always_comb begin // combinatorial arburst
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arburst = 2'bxx;
	arburst = _1;
end
always_comb begin // combinatorial arprot
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arprot = 3'bxxx;
	arprot = _2;
end
always_comb begin // combinatorial arcache
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arcache = 4'bxxxx;
	arcache = _3;
end
always_comb begin // combinatorial arqos
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arqos = 4'dx;
	arqos = 1'd0;
end
always_comb begin // combinatorial arlock
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arlock = 1'bx;
	arlock = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arlock = arlock;
end
always_comb begin // combinatorial arregion
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arregion = 4'dx;
	arregion = 1'd0;
end
always_comb begin // combinatorial rready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rready = 1'bx;
	rready = 1'b0;
	if(_13) rready = 1'b1;
	if(!_13) rready = do_read;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rready = rready;
end
always_comb begin // combinatorial _rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rresp = 2'bxx;
	_rresp = rresp;
end
always_comb begin // combinatorial _rlast
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_rlast = 1'bx;
	_rlast = rlast;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_rlast = _rlast;
end
always_comb begin // combinatorial fire
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	fire = 1'bx;
	if(request) fire = arready;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	fire = fire;
end
always_comb begin // combinatorial do_read
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	do_read = 1'bx;
	if(read) do_read = 1'b1;
	if(!read) do_read = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	do_read = do_read;
end
always_comb begin // combinatorial do_read_was_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	do_read_was_valid = 1'bx;
	if(_13) do_read_was_valid = 1'b0;
	if(!_13) do_read_was_valid = rvalid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	do_read_was_valid = do_read_was_valid;
end
always_comb begin // combinatorial do_read_data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	do_read_data = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(!_13) if(_25) do_read_data[_v0] = _27[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(!_13) if(_25) do_read_data[32 + _v0] = _28[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(!_13) if(_25) do_read_data[64 + _v0] = _29[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(!_13) if(_25) do_read_data[96 + _v0] = _30[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(!_13) if(_25) do_read_data[128 + _v0] = _31[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(!_13) if(_25) do_read_data[160 + _v0] = _32[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(!_13) if(_25) do_read_data[192 + _v0] = _33[_v0];
end
	for(int _v0 = 0; _v0 < 32; _v0 = _v0 + 1) begin
if(!_13) if(_25) do_read_data[224 + _v0] = rdata[_v0];
end
end
always_ff @(posedge aclk) begin // state stored_part_idx
	if(_13) if(rvalid) stored_part_idx <= _20;
	if(!_13) if(_25) stored_part_idx <= 1'd0;
	if(_36) stored_part_idx <= 1'd0;
end
always_ff @(posedge aclk) begin // state stored_parts
	if(_13) if(rvalid) stored_parts[idx] <= rdata;
end
always_comb begin // combinatorial idx
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	idx = 3'dx;
	if(_13) if(rvalid) idx = _IntNarrow_out;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 3'dx;
	if(_13) if(rvalid) _IntNarrow_in = stored_part_idx;
end
always_comb begin // combinatorial read_valid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	read_valid = 1'bx;
	if(read) read_valid = do_read_was_valid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	read_valid = read_valid;
end
always_comb begin // combinatorial data
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	data = '{32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx, 32'dx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(read) if(do_read_was_valid) data[_v0] = _FromBits_value[_v0];
end
end
always_comb begin // combinatorial _FromBits_bits
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_FromBits_bits = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(read) if(do_read_was_valid) _FromBits_bits = do_read_data;
end
endmodule

// FromBits #(T: type int #(FROM: 0, TO: 4294967296)[8])
module FromBits_T_type_int_FROM_0_TO_4294967296_8(
	input clk,
	input wire[255:0] bits,
	output /*mux_wire*/ logic[31:0] value[7:0]
);

genvar _g0;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign value[_g0] = bits[(_g0) * 32 +: 32];
end
endgenerate
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 8, FROM: 0, TO: 7)
module IntNarrow_FROM_I_0_TO_I_8_FROM_0_TO_7(
	input clk,
	input wire[2:0] in,
	output /*mux_wire*/ logic[2:0] out
);

	assign out = in;
endmodule

// axi_ctrl_slave #(NUM_INPUT_REGS: 8, NUM_OUTPUT_REGS: 1, ADDR_WIDTH: 12, AXI_WIDTH: 32)
module axi_ctrl_slave_NUM_INPUT_REGS_8_NUM_OUTPUT_REGS_1_ADDR_WIDTH_12_AXI_WIDTH_32(
	input aclk,
	input wire aresetn,
	input wire[11:0] awaddr,
	input wire awvalid,
	output /*mux_wire*/ logic awready,
	input wire[31:0] wdata,
	input wire[3:0] wstrb,
	input wire wvalid,
	output /*mux_wire*/ logic wready,
	output /*mux_wire*/ logic[1:0] bresp,
	output /*mux_wire*/ logic bvalid,
	input wire bready,
	input wire[11:0] araddr,
	input wire arvalid,
	output /*mux_wire*/ logic arready,
	output /*mux_wire*/ logic[31:0] rdata,
	output /*mux_wire*/ logic[1:0] rresp,
	output /*mux_wire*/ logic rvalid,
	input wire rready,
	output /*state*/ logic[31:0] input_regs[7:0],
	output /*mux_wire*/ logic start,
	input wire finish,
	input wire[31:0] output_regs[0:0]
);

genvar _g0;
/*state*/ logic[31:0] stored_output_regs[0:0];
/*state*/ logic reg_ctrl_ap_idle;
/*state*/ logic reg_ctrl_ap_done;
/*mux_wire*/ logic reg_ctrl_ap_ready;
/*state*/ logic reg_ctrl_ap_start;
/*state*/ logic[9:0] stored_addr;
/*state*/ logic stored_addr_valid;
/*state*/ logic[1:0] last_bresp;
/*state*/ logic last_werr_valid;
wire _4;
assign _4 = !stored_addr_valid;
wire _6;
assign _6 = _4 & aresetn;
wire _9;
assign _9 = !last_werr_valid;
wire _10;
assign _10 = stored_addr_valid & _9;
wire _15;
assign _15 = awready & awvalid;
wire[9:0] _17;
assign _17 = awaddr / 3'd4;
wire _20;
assign _20 = wready & wvalid;
localparam[1:0] RESP_SLVERR = 2'b10;
wire _22;
assign _22 = stored_addr == 1'd0;
wire _23 = wstrb[0];
wire _24 = wdata[0];
wire _25;
assign _25 = _23 & _24;
localparam[1:0] RESP_OKAY = 2'b00;
wire _28;
assign _28 = stored_addr >= 3'd4;
wire _31;
assign _31 = stored_addr < 4'd12;
wire _32;
assign _32 = _28 & _31;
/*mux_wire*/ logic[2:0] write_idx;
/*mux_wire*/ logic[9:0] _IntNarrow_in;
wire[3:0] _IntNarrow_out;
wire[2:0] _34;
assign _34 = _IntNarrow_out - 3'd4;
wire _35 = wstrb[0];
wire[7:0] _37;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _37[_g0] = wdata[_g0];
end
endgenerate
wire _38 = wstrb[1];
wire[7:0] _40;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _40[_g0] = wdata[8 + _g0];
end
endgenerate
wire _41 = wstrb[2];
wire[7:0] _43;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _43[_g0] = wdata[16 + _g0];
end
endgenerate
wire _44 = wstrb[3];
wire[7:0] _46;
generate
for(_g0 = 0; _g0 < 8; _g0 = _g0 + 1) begin
assign _46[_g0] = wdata[24 + _g0];
end
endgenerate
localparam[1:0] RESP_OKAY_2 = 2'b00;
wire _49;
assign _49 = bready & bvalid;
/*state*/ logic last_rdata_valid;
/*state*/ logic[31:0] last_rdata;
/*state*/ logic[1:0] last_rresp;
/*mux_wire*/ logic[31:0] regs_read_multiplexer[8:0];
wire _55;
assign _55 = !last_rdata_valid;
wire _57;
assign _57 = _55 & aresetn;
wire _61;
assign _61 = arready & arvalid;
localparam[1:0] RESP_SLVERR_2 = 2'b10;
/*mux_wire*/ logic[9:0] read_addr;
wire[9:0] _63;
assign _63 = araddr / 3'd4;
wire _65;
assign _65 = read_addr == 1'd0;
/*mux_wire*/ logic _Repeat_v;
wire[27:0] _Repeat_result;
localparam[1:0] RESP_OKAY_3 = 2'b00;
wire _72;
assign _72 = read_addr >= 3'd4;
wire _75;
assign _75 = read_addr < 4'd13;
wire _76;
assign _76 = _72 & _75;
/*mux_wire*/ logic[3:0] read_idx;
/*mux_wire*/ logic[9:0] _IntNarrow_2_in;
wire[3:0] _IntNarrow_2_out;
wire[3:0] _78;
assign _78 = _IntNarrow_2_out - 3'd4;
wire[31:0] _80 = regs_read_multiplexer[read_idx];
localparam[1:0] RESP_OKAY_4 = 2'b00;
wire _83;
assign _83 = rready & rvalid;
/*mux_wire*/ logic _cross_finish_in;
/*mux_wire*/ logic[31:0] _cross_finish_data_in[0:0];
wire _cross_finish_out;
wire[31:0] _cross_finish_data_out[0:0];
/*mux_wire*/ logic[31:0] output_regs_vs[0:0];
wire _89;
assign _89 = !aresetn;
/*mux_wire*/ logic _Repeat_2_v;
wire[31:0] _Repeat_2_result;
/*mux_wire*/ logic[31:0] _Repeat_3_v;
wire[31:0] _Repeat_3_result[7:0];
/*mux_wire*/ logic _Repeat_4_v;
wire[31:0] _Repeat_4_result;
/*mux_wire*/ logic[31:0] _Repeat_5_v;
wire[31:0] _Repeat_5_result[0:0];
IntNarrow_FROM_I_0_TO_I_1024_FROM_4_TO_12 IntNarrow(
	.clk(aclk),
	.in(_IntNarrow_in),
	.out(_IntNarrow_out)
);
Repeat_T_type_bool_SIZE_28 Repeat(
	.clk(aclk),
	.v(_Repeat_v),
	.result(_Repeat_result)
);
IntNarrow_FROM_I_0_TO_I_1024_FROM_4_TO_13 IntNarrow_2(
	.clk(aclk),
	.in(_IntNarrow_2_in),
	.out(_IntNarrow_2_out)
);
CrossAction_T_type_bool_32_1 cross_finish(
	.in_clk(aclk),
	.in(_cross_finish_in),
	.data_in(_cross_finish_data_in),
	.out(_cross_finish_out),
	.data_out(_cross_finish_data_out)
);
Repeat_T_type_bool_SIZE_32 Repeat_2(
	.clk(aclk),
	.v(_Repeat_2_v),
	.result(_Repeat_2_result)
);
Repeat_T_type_bool_32_SIZE_8 Repeat_3(
	.clk(aclk),
	.v(_Repeat_3_v),
	.result(_Repeat_3_result)
);
Repeat_T_type_bool_SIZE_32 Repeat_4(
	.clk(aclk),
	.v(_Repeat_4_v),
	.result(_Repeat_4_result)
);
Repeat_T_type_bool_32_SIZE_1 Repeat_5(
	.clk(aclk),
	.v(_Repeat_5_v),
	.result(_Repeat_5_result)
);
always_comb begin // combinatorial awready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	awready = 1'bx;
	awready = 1'b0;
	awready = _6;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	awready = awready;
end
always_comb begin // combinatorial wready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	wready = 1'bx;
	wready = 1'b0;
	wready = _10;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	wready = wready;
end
always_comb begin // combinatorial bresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	bresp = 2'bxx;
	bresp = last_bresp;
end
always_comb begin // combinatorial bvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	bvalid = 1'bx;
	bvalid = 1'b0;
	bvalid = last_werr_valid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	bvalid = bvalid;
end
always_comb begin // combinatorial arready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	arready = 1'bx;
	arready = 1'b0;
	arready = _57;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	arready = arready;
end
always_comb begin // combinatorial rdata
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rdata = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	rdata = last_rdata;
end
always_comb begin // combinatorial rresp
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rresp = 2'bxx;
	rresp = last_rresp;
end
always_comb begin // combinatorial rvalid
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	rvalid = 1'bx;
	rvalid = 1'b0;
	rvalid = last_rdata_valid;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	rvalid = rvalid;
end
always_ff @(posedge aclk) begin // state stored_output_regs
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_cross_finish_out) stored_output_regs[_v0] <= output_regs_vs[_v0];
end
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_89) stored_output_regs[_v0] <= _Repeat_5_result[_v0];
end
end
always_ff @(posedge aclk) begin // state input_regs
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_20) if(_32) if(_35) input_regs[write_idx][_v0] <= _37[_v0];
end
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_20) if(_32) if(_38) input_regs[write_idx][8 + _v0] <= _40[_v0];
end
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_20) if(_32) if(_41) input_regs[write_idx][16 + _v0] <= _43[_v0];
end
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_20) if(_32) if(_44) input_regs[write_idx][24 + _v0] <= _46[_v0];
end
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
if(_89) input_regs[_v0] <= _Repeat_3_result[_v0];
end
end
always_comb begin // combinatorial start
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	start = 1'bx;
	start = 1'b0;
	if(_20) if(_22) if(_25) start = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	start = start;
end
always_ff @(posedge aclk) begin // state reg_ctrl_ap_idle
	if(_20) if(_22) if(_25) reg_ctrl_ap_idle <= 1'b0;
	if(_61) if(_65) if(reg_ctrl_ap_done) reg_ctrl_ap_idle <= 1'b1;
	if(_cross_finish_out) reg_ctrl_ap_idle <= 1'b0;
	if(_89) reg_ctrl_ap_idle <= 1'b1;
end
always_ff @(posedge aclk) begin // state reg_ctrl_ap_done
	if(_61) if(_65) reg_ctrl_ap_done <= 1'b0;
	if(_cross_finish_out) reg_ctrl_ap_done <= 1'b1;
	if(_89) reg_ctrl_ap_done <= 1'b0;
end
always_comb begin // combinatorial reg_ctrl_ap_ready
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	reg_ctrl_ap_ready = 1'bx;
	reg_ctrl_ap_ready = reg_ctrl_ap_done;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	reg_ctrl_ap_ready = reg_ctrl_ap_ready;
end
always_ff @(posedge aclk) begin // state reg_ctrl_ap_start
	if(_20) if(_22) if(_25) reg_ctrl_ap_start <= 1'b1;
	if(_cross_finish_out) reg_ctrl_ap_start <= 1'b0;
	if(_89) reg_ctrl_ap_start <= 1'b0;
end
always_ff @(posedge aclk) begin // state stored_addr
	if(_15) stored_addr <= _17;
end
always_ff @(posedge aclk) begin // state stored_addr_valid
	if(_15) stored_addr_valid <= 1'b1;
	if(_20) stored_addr_valid <= 1'b0;
	if(_89) stored_addr_valid <= 1'b0;
end
always_ff @(posedge aclk) begin // state last_bresp
	if(_20) last_bresp <= RESP_SLVERR;
	if(_20) if(_22) last_bresp <= RESP_OKAY;
	if(_20) if(_32) last_bresp <= RESP_OKAY_2;
end
always_ff @(posedge aclk) begin // state last_werr_valid
	if(_20) last_werr_valid <= 1'b1;
	if(_49) last_werr_valid <= 1'b0;
	if(_89) last_werr_valid <= 1'b0;
end
always_comb begin // combinatorial write_idx
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	write_idx = 3'dx;
	if(_20) if(_32) write_idx = _34;
end
always_comb begin // combinatorial _IntNarrow_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_in = 10'dx;
	if(_20) if(_32) _IntNarrow_in = stored_addr;
end
always_ff @(posedge aclk) begin // state last_rdata_valid
	if(_61) last_rdata_valid <= 1'b1;
	if(_83) last_rdata_valid <= 1'b0;
	if(_89) last_rdata_valid <= 1'b0;
end
always_ff @(posedge aclk) begin // state last_rdata
	if(_61) if(_65) last_rdata[0] <= reg_ctrl_ap_start;
	if(_61) if(_65) last_rdata[1] <= reg_ctrl_ap_done;
	if(_61) if(_65) last_rdata[2] <= reg_ctrl_ap_idle;
	if(_61) if(_65) last_rdata[3] <= reg_ctrl_ap_ready;
	for(int _v0 = 0; _v0 < 28; _v0 = _v0 + 1) begin
if(_61) if(_65) last_rdata[4 + _v0] <= _Repeat_result[_v0];
end
	if(_61) if(_76) last_rdata <= _80;
end
always_ff @(posedge aclk) begin // state last_rresp
	if(_61) last_rresp <= RESP_SLVERR_2;
	if(_61) if(_65) last_rresp <= RESP_OKAY_3;
	if(_61) if(_76) last_rresp <= RESP_OKAY_4;
end
always_comb begin // combinatorial regs_read_multiplexer
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	regs_read_multiplexer = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 8; _v0 = _v0 + 1) begin
regs_read_multiplexer[_v0] = input_regs[_v0];
end
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
regs_read_multiplexer[8 + _v0] = stored_output_regs[_v0];
end
end
always_comb begin // combinatorial read_addr
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	read_addr = 10'dx;
	if(_61) read_addr = _63;
end
always_comb begin // combinatorial _Repeat_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_v = 1'bx;
	if(_61) if(_65) _Repeat_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_v = _Repeat_v;
end
always_comb begin // combinatorial read_idx
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	read_idx = 4'dx;
	if(_61) if(_76) read_idx = _78;
end
always_comb begin // combinatorial _IntNarrow_2_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_IntNarrow_2_in = 10'dx;
	if(_61) if(_76) _IntNarrow_2_in = read_addr;
end
always_comb begin // combinatorial _cross_finish_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_finish_in = 1'bx;
	_cross_finish_in = 1'b0;
	if(finish) _cross_finish_in = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_finish_in = _cross_finish_in;
end
always_comb begin // combinatorial _cross_finish_data_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_finish_data_in = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(finish) _cross_finish_data_in[_v0] = output_regs[_v0];
end
end
always_comb begin // combinatorial output_regs_vs
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	output_regs_vs = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_cross_finish_out) output_regs_vs[_v0] = _cross_finish_data_out[_v0];
end
end
always_comb begin // combinatorial _Repeat_2_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_2_v = 1'bx;
	if(_89) _Repeat_2_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_2_v = _Repeat_2_v;
end
always_comb begin // combinatorial _Repeat_3_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_3_v = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_89) _Repeat_3_v = _Repeat_2_result;
end
always_comb begin // combinatorial _Repeat_4_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_4_v = 1'bx;
	if(_89) _Repeat_4_v = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_Repeat_4_v = _Repeat_4_v;
end
always_comb begin // combinatorial _Repeat_5_v
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_Repeat_5_v = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	if(_89) _Repeat_5_v = _Repeat_4_result;
end
endmodule

// Repeat #(T: type bool #()[32], SIZE: 1)
module Repeat_T_type_bool_32_SIZE_1(
	input clk,
	input wire[31:0] v,
	output /*mux_wire*/ logic[31:0] result[0:0]
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	result[0] = v;
end
endmodule

// Repeat #(T: type bool #()[32], SIZE: 8)
module Repeat_T_type_bool_32_SIZE_8(
	input clk,
	input wire[31:0] v,
	output /*mux_wire*/ logic[31:0] result[7:0]
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx, 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
	result[4] = v;
	result[5] = v;
	result[6] = v;
	result[7] = v;
end
endmodule

// Repeat #(T: type bool #(), SIZE: 32)
module Repeat_T_type_bool_SIZE_32(
	input clk,
	input wire v,
	output /*mux_wire*/ logic[31:0] result
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
	result[4] = v;
	result[5] = v;
	result[6] = v;
	result[7] = v;
	result[8] = v;
	result[9] = v;
	result[10] = v;
	result[11] = v;
	result[12] = v;
	result[13] = v;
	result[14] = v;
	result[15] = v;
	result[16] = v;
	result[17] = v;
	result[18] = v;
	result[19] = v;
	result[20] = v;
	result[21] = v;
	result[22] = v;
	result[23] = v;
	result[24] = v;
	result[25] = v;
	result[26] = v;
	result[27] = v;
	result[28] = v;
	result[29] = v;
	result[30] = v;
	result[31] = v;
end
endmodule

// CrossAction #(T: type bool #()[32][1])
module CrossAction_T_type_bool_32_1(
	input in_clk,
	input wire in,
	input wire[31:0] data_in[0:0],
	output /*mux_wire*/ logic out,
	output /*mux_wire*/ logic[31:0] data_out[0:0]
);

/*mux_wire*/ logic _cross_valid_in;
/*mux_wire*/ logic[31:0] _cross_data_in[0:0];
wire _cross_valid_out;
wire[31:0] _cross_data_out[0:0];
CrossDomain_T_type_bool cross_valid(
	.in_clk(in_clk),
	.in(_cross_valid_in),
	.out(_cross_valid_out)
);
CrossDomain_T_type_bool_32_1 cross_data(
	.in_clk(in_clk),
	.in(_cross_data_in),
	.out(_cross_data_out)
);
always_comb begin // combinatorial _cross_valid_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_valid_in = 1'bx;
	if(in) _cross_valid_in = 1'b1;
	if(!in) _cross_valid_in = 1'b0;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	_cross_valid_in = _cross_valid_in;
end
always_comb begin // combinatorial _cross_data_in
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	_cross_data_in = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(in) _cross_data_in[_v0] = data_in[_v0];
end
end
always_comb begin // combinatorial out
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	out = 1'bx;
	out = 1'b0;
	if(_cross_valid_out) out = 1'b1;
	// PATCH Vivado 23.1 Simulator Bug: 1-bit Conditional Assigns become don't care
	out = out;
end
always_comb begin // combinatorial data_out
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	data_out = '{32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx};
	for(int _v0 = 0; _v0 < 1; _v0 = _v0 + 1) begin
if(_cross_valid_out) data_out[_v0] = _cross_data_out[_v0];
end
end
endmodule

// CrossDomain #(T: type bool #()[32][1])
module CrossDomain_T_type_bool_32_1(
	input in_clk,
	input wire[31:0] in[0:0],
	output /*mux_wire*/ logic[31:0] out[0:0]
);

	assign out = in;
endmodule

// CrossDomain #(T: type bool #())
module CrossDomain_T_type_bool(
	input in_clk,
	input wire in,
	output /*mux_wire*/ logic out
);

	assign out = in;
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 1024, FROM: 4, TO: 13)
module IntNarrow_FROM_I_0_TO_I_1024_FROM_4_TO_13(
	input clk,
	input wire[9:0] in,
	output /*mux_wire*/ logic[3:0] out
);

	assign out = in;
endmodule

// Repeat #(T: type bool #(), SIZE: 28)
module Repeat_T_type_bool_SIZE_28(
	input clk,
	input wire v,
	output /*mux_wire*/ logic[27:0] result
);

always_comb begin // combinatorial result
	// Combinatorial wires are not defined when not valid. This is just so that the synthesis tool doesn't generate latches
	result = 28'bxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	result[0] = v;
	result[1] = v;
	result[2] = v;
	result[3] = v;
	result[4] = v;
	result[5] = v;
	result[6] = v;
	result[7] = v;
	result[8] = v;
	result[9] = v;
	result[10] = v;
	result[11] = v;
	result[12] = v;
	result[13] = v;
	result[14] = v;
	result[15] = v;
	result[16] = v;
	result[17] = v;
	result[18] = v;
	result[19] = v;
	result[20] = v;
	result[21] = v;
	result[22] = v;
	result[23] = v;
	result[24] = v;
	result[25] = v;
	result[26] = v;
	result[27] = v;
end
endmodule

// IntNarrow #(FROM_I: 0, TO_I: 1024, FROM: 4, TO: 12)
module IntNarrow_FROM_I_0_TO_I_1024_FROM_4_TO_12(
	input clk,
	input wire[9:0] in,
	output /*mux_wire*/ logic[3:0] out
);

	assign out = in;
endmodule

